current-steering dac inl test

*.option gmin=1e-19 reltol=200u abstol=100f vntol=100n seed=2

.param mc_mm_switch = 1
.param vdd = 1.5

vdd vdd 0 dc vdd
xdac1 vdd 0 b16 b15 b14 b13 b12 b11 bb16 bb15 bb14 bb13 bb12 bb11 outp1 outn1 dac
xdac2 vdd 0 b26 b25 b24 b23 b22 b21 bb26 bb25 bb24 bb23 bb22 bb21 outp2 outn2 dac
rlp1 outp1 0 0.02
rln1 outn1 0 0.02
rlp2 outp2 0 0.02
rln2 outn2 0 0.02
e1 out1 0 outp1 outn1 10
rl1 out1 0 1k
e2 out2 0 outp2 outn2 10
rl2 out 0 1k

.subckt pfet d g s b
.param mfac = 1
xm d g s b sky130_fd_pr__pfet_01v8_lvt l=350n w=550n as=145.75f ad=145.75f ps=1.63u pd=1.63u mult=mfac m=mfac
.ends

.subckt cell vdd vss bp b bb outp outn weight=1
c1 d1 vdd '20f*weight'
c2 bp vdd '20f*weight'
xm1 d1 bp vdd vdd pfet mfac=weight
xm2p outp bb d1 vdd pfet mfac=weight
xm2n outn b d1 vdd pfet mfac=weight
.ends

.subckt dac vdd vss b6 b5 b4 b3 b2 b1 bb6 bb5 bb4 bb3 bb2 bb1 outp outn
xmb1 bp bp vdd vdd pfet mfac=1
xmb2 0 0 bp vdd pfet mfac=1
xdc1 vdd 0 bp b1 bb1 outp outn cell weight=1
xdc2 vdd 0 bp b2 bb2 outp outn cell weight=2
xdc3 vdd 0 bp b3 bb3 outp outn cell weight=4
xdc4 vdd 0 bp b4 bb4 outp outn cell weight=8
xdc5 vdd 0 bp b5 bb5 outp outn cell weight=16
xdc6 vdd 0 bp b6 bb6 outp outn cell weight=32
.ends

.param
+ sky130_fd_pr__pfet_01v8_lvt__ajunction_mult = 9.9626e-1
+ sky130_fd_pr__pfet_01v8_lvt__pjunction_mult = 1.0009e+0
+ sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff = .73e-6
+ sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__wlod_diff = .0e-6
+ sky130_fd_pr__pfet_01v8_lvt__ku0_diff = 5.9e-8
+ sky130_fd_pr__pfet_01v8_lvt__lku0_diff = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__wku0_diff = 0.0
+ sky130_fd_pr__pfet_01v8_lvt__kvsat_diff = .0e-6
+ sky130_fd_pr__pfet_01v8_lvt__kvth0_diff = 1.76e-8

.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope=3.689e-09
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope1=1.489e-08
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope2=1.689e-08
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope3=2.389e-08
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope=1.389e-08
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope1=9.789e-09
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope2=1.089e-08
.param sky130_fd_pr__pfet_01v8_lvt__lint_slope=0
.param sky130_fd_pr__pfet_01v8_lvt__wint_slope=0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope=0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope=0.0

.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre = 0.0

.subckt  sky130_fd_pr__pfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1
msky130_fd_pr__pfet_01v8_lvt d g s b sky130_fd_pr__pfet_01v8_lvt__model l = {l} w = {w} nf = {nf} ad = {ad} as = {as} pd = {pd} ps = {ps} nrd = {nrd} nrs = {nrs} sa = {sa} sb = {sb} sd = {sd}
.model sky130_fd_pr__pfet_01v8_lvt__model pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 2.8e-9
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 7.476e-9
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre)
+ toxe = {4.23e-09+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(4.23e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(l*w*mult)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre)
+ vth0 = {-1.782289999e-01+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(l*w*mult))} lvth0 = -7.222604304e-08 wvth0 = -1.348985490e-07 pvth0 = 4.954643417e-14
+ k1 = 0.64774
+ k2 = -4.695523411e-02 lk2 = 4.071953082e-09 wk2 = -1.048260450e-08 pk2 = 6.073815561e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.729186447e+05 lvsat = -1.976658997e-02 wvsat = -6.300395056e-02 pvsat = 1.733533569e-8
+ ua = -3.076683126e-09 lua = 6.229870963e-17 wua = 2.386014056e-16 pua = -1.060940094e-22
+ ub = 2.612994519e-18 lub = 1.905974519e-25 wub = -8.036427329e-26 pub = 6.115694775e-32
+ uc = 1.607392219e-11 luc = 1.380586924e-17 wuc = 4.015260322e-17 puc = -1.359944388e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 9.335311068e-04 lu0 = 6.553868693e-10 wu0 = 1.170785149e-09 pu0 = -4.005819962e-16
+ a0 = 1.1627
+ keta = -1.727227166e-02 lketa = 1.876040360e-09 wketa = 2.914551807e-09 pketa = -1.003771642e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -7.446080985e-01 lags = 3.523067795e-07 wags = 9.865926523e-07 pags = -3.470390885e-13
+ b0 = 7.894683512e-07 lb0 = -4.041704517e-13 wb0 = -7.386199123e-13 pb0 = 3.251555372e-19
+ b1 = -1.841702328e-06 lb1 = 7.894705525e-13 wb1 = 1.711615945e-12 pb1 = -6.725137054e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre)
+ voff = {-0.1819+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(l*w*mult))}
*(mismatch parameter sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre)
+ nfactor = {2.5373+MC_MM_SWITCH*AGAUSS(0,1.0,1)*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(l*w*mult))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.703778191e-03 lpdiblc2 = 9.640935270e-09 wpdiblc2 = -4.489995143e-08 ppdiblc2 = 3.814731091e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.509909476e-01 ldelta = -2.800512739e-08 wdelta = -6.545113965e-08 pdelta = 1.652434138e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.924373247e-01 lkt1 = 6.087865133e-08 wkt1 = 1.276072598e-07 pkt1 = -4.798161401e-14
+ kt2 = 1.626020472e-01 lkt2 = -8.539089664e-08 wkt2 = -1.326603614e-07 pkt2 = 4.568822846e-14
+ at = -4.433949910e+04 lat = 2.869593405e-02 wat = 1.874991537e-01 pat = -6.980799686e-8
+ ute = -8.127409949e-01 lute = 2.067746586e-07 wute = 5.193692717e-07 pute = -1.788707772e-13
+ ua1 = 1.972651465e-09 lua1 = -4.303214166e-16 wua1 = -6.685325589e-16 pua1 = 2.302426133e-22
+ ub1 = -2.955731024e-18 lub1 = 9.378910967e-25 wub1 = 1.375089403e-24 pub1 = -4.735807904e-31
+ uc1 = -1.642735167e-10 luc1 = 6.690779914e-17 wuc1 = 1.039456565e-16 puc1 = -3.579888411e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 2.0e-11
+ cgso = 2.0e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = -1.2e-8
+ dwc = 0.0
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007653568198
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 9.1602368e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.39155046e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8_lvt


.option method=trap TRTOL=5 gmin=1e-19 reltol=200u abstol=100f vntol=100n seed=2

.control
tran 10u 0.006999186686686687
write $inputdir/cs_dac_06bit_2ch_TRAN_ngspice_batch.bin v(out1) v(out2)
.endc

vb11 b11 0 pwl 0,0  0.9770400400400401u,0 0.97804004004004u,1.5 1.95458008008008u,1.5 1.95558008008008u,0 2.93212012012012u,0 2.9331201201201202u,1.5 3.90966016016016u,1.5 3.9106601601601603u,0 4.8872002002002u,0 4.8882002002002u,1.5 9.7749004004004u,1.5 9.7759004004004u,0 11.72998048048048u,0 11.730980480480481u,1.5 12.70752052052052u,1.5 12.708520520520521u,0 13.68506056056056u,0 13.686060560560561u,1.5 17.59522072072072u,1.5 17.59622072072072u,0 18.572760760760765u,0 18.573760760760763u,1.5 25.415541041041042u,1.5 25.41654104104104u,0 26.393081081081085u,0 26.394081081081083u,1.5 27.370621121121122u,1.5 27.37162112112112u,0 28.348161161161162u,0 28.34916116116116u,1.5 30.303241241241246u,1.5 30.304241241241243u,0 31.280781281281282u,0 31.28178128128128u,1.5 33.23586136136136u,1.5 33.23686136136136u,0 35.19094144144144u,0 35.19194144144144u,1.5 36.16848148148148u,1.5 36.16948148148148u,0 37.146021521521526u,0 37.14702152152153u,1.5 39.1011016016016u,1.5 39.1021016016016u,0 40.07864164164164u,0 40.07964164164164u,1.5 42.03372172172172u,1.5 42.03472172172172u,0 44.966341841841846u,0 44.96734184184185u,1.5 45.94388188188188u,1.5 45.944881881881884u,0 47.89896196196196u,0 47.899961961961964u,1.5 48.876502002002u,1.5 48.877502002002004u,0 50.83158208208208u,0 50.832582082082084u,1.5 52.786662162162166u,1.5 52.78766216216217u,0 53.7642022022022u,0 53.765202202202204u,1.5 54.74174224224224u,1.5 54.742742242242244u,0 55.71928228228228u,0 55.720282282282284u,1.5 58.6519024024024u,1.5 58.652902402402404u,0 59.62944244244244u,0 59.630442442442444u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 71.35992292292292u,0 71.36092292292292u,1.5 72.33746296296296u,1.5 72.33846296296296u,0 76.24762312312312u,0 76.24862312312312u,1.5 78.2027032032032u,1.5 78.2037032032032u,0 80.15778328328328u,0 80.15878328328328u,1.5 85.04548348348348u,1.5 85.04648348348348u,0 86.02302352352352u,0 86.02402352352352u,1.5 87.00056356356356u,1.5 87.00156356356356u,0 90.91072372372372u,0 90.91172372372372u,1.5 92.8658038038038u,1.5 92.8668038038038u,0 94.82088388388388u,0 94.82188388388388u,1.5 95.79842392392392u,1.5 95.79942392392392u,0 96.77596396396396u,0 96.77696396396396u,1.5 97.753504004004u,1.5 97.754504004004u,0 98.73104404404404u,0 98.73204404404404u,1.5 100.68612412412412u,1.5 100.68712412412413u,0 101.66366416416416u,0 101.66466416416417u,1.5 104.59628428428428u,1.5 104.59728428428429u,0 106.55136436436436u,0 106.55236436436437u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 109.48398448448448u,0 109.48498448448449u,1.5 111.43906456456456u,1.5 111.44006456456457u,0 114.37168468468468u,0 114.37268468468469u,1.5 115.34922472472472u,1.5 115.35022472472473u,0 117.3043048048048u,0 117.3053048048048u,1.5 123.16954504504503u,1.5 123.17054504504503u,0 124.14708508508508u,0 124.14808508508509u,1.5 125.12462512512512u,1.5 125.12562512512513u,0 127.07970520520522u,0 127.08070520520522u,1.5 128.05724524524524u,1.5 128.05824524524522u,0 130.01232532532532u,0 130.0133253253253u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 136.85510560560562u,0 136.8561056056056u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 139.78772572572572u,0 139.7887257257257u,1.5 140.76526576576578u,1.5 140.76626576576575u,0 141.74280580580583u,0 141.7438058058058u,1.5 142.72034584584586u,1.5 142.72134584584583u,0 143.69788588588588u,0 143.69888588588586u,1.5 144.67542592592594u,1.5 144.6764259259259u,0 145.65296596596596u,0 145.65396596596594u,1.5 150.54066616616618u,1.5 150.54166616616615u,0 152.49574624624626u,0 152.49674624624623u,1.5 153.4732862862863u,1.5 153.4742862862863u,0 156.40590640640642u,0 156.4069064064064u,1.5 158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 165.20376676676676u,1.5 165.20476676676674u,0 168.1363868868869u,0 168.13738688688687u,1.5 169.11392692692695u,1.5 169.11492692692693u,0 170.09146696696698u,0 170.09246696696695u,1.5 174.97916716716716u,1.5 174.98016716716714u,0 178.88932732732735u,0 178.89032732732733u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 185.73210760760762u,0 185.7331076076076u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 189.64226776776778u,1.5 189.64326776776775u,0 190.6198078078078u,0 190.62080780780778u,1.5 191.59734784784786u,1.5 191.59834784784783u,0 192.57488788788788u,0 192.57588788788786u,1.5 194.529967967968u,1.5 194.53096796796797u,0 197.4625880880881u,0 197.46358808808807u,1.5 198.44012812812815u,1.5 198.44112812812813u,0 201.37274824824826u,0 201.37374824824823u,1.5 203.32782832832834u,1.5 203.3288283283283u,0 204.3053683683684u,0 204.30636836836837u,1.5 207.2379884884885u,1.5 207.23898848848847u,0 208.21552852852852u,0 208.2165285285285u,1.5 210.17060860860863u,1.5 210.1716086086086u,0 211.1481486486487u,0 211.14914864864866u,1.5 212.12568868868868u,1.5 212.12668868868866u,0 214.0807687687688u,0 214.08176876876877u,1.5 218.96846896896898u,1.5 218.96946896896895u,0 219.94600900900903u,0 219.947009009009u,1.5 220.92354904904906u,1.5 220.92454904904903u,0 223.85616916916916u,0 223.85716916916914u,1.5 229.72140940940943u,1.5 229.7224094094094u,0 230.69894944944946u,0 230.69994944944943u,1.5 231.6764894894895u,1.5 231.6774894894895u,0 233.63156956956956u,0 233.63256956956954u,1.5 234.60910960960962u,1.5 234.6101096096096u,0 236.5641896896897u,0 236.56518968968967u,1.5 237.54172972972972u,1.5 237.5427297297297u,0 238.51926976976978u,0 238.52026976976975u,1.5 239.4968098098098u,1.5 239.49780980980978u,0 240.47434984984986u,0 240.47534984984983u,1.5 241.4518898898899u,1.5 241.4528898898899u,0 242.42942992992997u,0 242.43042992992994u,1.5 243.40696996996996u,1.5 243.40796996996994u,0 245.36205005005007u,0 245.36305005005005u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 256.11499049049047u,0 256.11599049049045u,1.5 259.04761061061066u,1.5 259.04861061061064u,0 260.02515065065063u,0 260.0261506506506u,1.5 261.00269069069066u,1.5 261.00369069069063u,0 261.98023073073074u,0 261.9812307307307u,1.5 263.93531081081085u,1.5 263.9363108108108u,0 265.8903908908909u,0 265.8913908908909u,1.5 270.77809109109114u,1.5 270.7790910910911u,0 271.75563113113117u,0 271.75663113113114u,1.5 272.73317117117114u,1.5 272.7341711711711u,0 275.6657912912913u,0 275.6667912912913u,1.5 279.57595145145143u,1.5 279.5769514514514u,0 280.5534914914915u,0 280.5544914914915u,1.5 281.53103153153154u,1.5 281.5320315315315u,0 282.50857157157157u,0 282.50957157157154u,1.5 283.48611161161165u,1.5 283.4871116116116u,0 287.39627177177175u,0 287.3972717717717u,1.5 289.35135185185186u,1.5 289.35235185185184u,0 290.32889189189194u,0 290.3298918918919u,1.5 294.23905205205205u,1.5 294.240052052052u,0 297.17167217217224u,0 297.1726721721722u,1.5 298.1492122122122u,1.5 298.1502122122122u,0 300.1042922922923u,0 300.1052922922923u,1.5 302.0593723723724u,1.5 302.0603723723724u,0 304.0144524524524u,0 304.0154524524524u,1.5 307.92461261261263u,1.5 307.9256126126126u,0 308.90215265265266u,0 308.90315265265264u,1.5 313.78985285285285u,1.5 313.7908528528528u,0 314.76739289289293u,0 314.7683928928929u,1.5 315.74493293293295u,1.5 315.74593293293293u,0 317.700013013013u,0 317.701013013013u,1.5 318.67755305305303u,1.5 318.678553053053u,0 320.63263313313314u,0 320.6336331331331u,1.5 321.6101731731732u,1.5 321.6111731731732u,0 322.5877132132132u,0 322.58871321321317u,1.5 323.5652532532532u,1.5 323.5662532532532u,0 324.5427932932933u,0 324.5437932932933u,1.5 326.4978733733734u,1.5 326.4988733733734u,0 328.45295345345346u,0 328.45395345345344u,1.5 330.4080335335335u,1.5 330.4090335335335u,0 332.3631136136136u,0 332.3641136136136u,1.5 333.3406536536537u,1.5 333.3416536536537u,0 334.31819369369373u,0 334.3191936936937u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 336.2732737737738u,0 336.27427377377376u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 338.2283538538539u,0 338.22935385385387u,1.5 340.18343393393394u,1.5 340.1844339339339u,0 343.1160540540541u,0 343.11705405405405u,1.5 344.0935940940941u,1.5 344.0945940940941u,0 345.0711341341341u,0 345.0721341341341u,1.5 349.9588343343343u,1.5 349.9598343343343u,0 350.9363743743744u,0 350.9373743743744u,1.5 353.8689944944945u,1.5 353.86999449449445u,0 354.8465345345345u,0 354.8475345345345u,1.5 355.8240745745746u,1.5 355.82507457457456u,0 357.7791546546547u,0 357.78015465465467u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 367.55455505505506u,0 367.55555505505504u,1.5 368.5320950950951u,1.5 368.53309509509506u,0 371.4647152152152u,0 371.4657152152152u,1.5 372.44225525525525u,1.5 372.4432552552552u,0 375.3748753753754u,0 375.37587537537536u,1.5 378.3074954954955u,1.5 378.3084954954955u,0 380.26257557557557u,0 380.26357557557554u,1.5 381.2401156156156u,1.5 381.24111561561557u,0 386.1278158158158u,0 386.12881581581576u,1.5 388.0828958958959u,1.5 388.08389589589586u,0 390.037975975976u,0 390.038975975976u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 395.90321621621626u,1.5 395.90421621621624u,0 396.8807562562563u,0 396.88175625625627u,1.5 398.83583633633634u,1.5 398.8368363363363u,0 399.81337637637637u,0 399.81437637637634u,1.5 400.79091641641645u,1.5 400.7919164164164u,0 401.7684564564565u,0 401.76945645645645u,1.5 402.7459964964965u,1.5 402.7469964964965u,0 403.7235365365366u,0 403.72453653653656u,1.5 404.70107657657655u,1.5 404.70207657657653u,0 406.65615665665666u,0 406.65715665665664u,1.5 407.6336966966967u,1.5 407.63469669669666u,0 409.5887767767768u,0 409.5897767767768u,1.5 410.5663168168168u,1.5 410.5673168168168u,0 411.54385685685685u,0 411.5448568568568u,1.5 412.5213968968969u,1.5 412.52239689689685u,0 414.476476976977u,0 414.47747697697696u,1.5 415.45401701701707u,1.5 415.45501701701704u,0 417.40909709709706u,0 417.41009709709704u,1.5 418.38663713713714u,1.5 418.3876371371371u,0 422.29679729729736u,0 422.29779729729734u,1.5 424.25187737737735u,1.5 424.25287737737733u,0 425.22941741741744u,0 425.2304174174174u,1.5 427.18449749749755u,1.5 427.1854974974975u,0 428.16203753753757u,0 428.16303753753755u,1.5 432.07219769769773u,1.5 432.0731976976977u,0 433.04973773773776u,0 433.05073773773773u,1.5 434.0272777777778u,1.5 434.02827777777776u,0 435.00481781781787u,0 435.00581781781784u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 437.93743793793794u,0 437.9384379379379u,1.5 438.91497797797797u,1.5 438.91597797797795u,0 449.6679184184184u,0 449.6689184184184u,1.5 450.64545845845845u,1.5 450.6464584584584u,0 451.62299849849853u,0 451.6239984984985u,1.5 452.60053853853856u,1.5 452.60153853853853u,0 453.5780785785786u,0 453.57907857857856u,1.5 455.53315865865864u,1.5 455.5341586586586u,0 456.5106986986987u,0 456.5116986986987u,1.5 460.4208588588588u,1.5 460.4218588588588u,0 461.3983988988989u,0 461.3993988988989u,1.5 462.37593893893893u,1.5 462.3769389389389u,0 463.353478978979u,0 463.354478978979u,1.5 466.28609909909915u,1.5 466.2870990990991u,0 468.2411791791792u,0 468.2421791791792u,1.5 470.19625925925925u,1.5 470.1972592592592u,0 471.17379929929933u,0 471.1747992992993u,1.5 472.15133933933936u,1.5 472.15233933933933u,0 474.1064194194194u,0 474.1074194194194u,1.5 475.08395945945944u,1.5 475.0849594594594u,0 476.0614994994995u,0 476.0624994994995u,1.5 478.0165795795796u,1.5 478.0175795795796u,0 484.8593598598599u,0 484.8603598598599u,1.5 485.8368998998999u,1.5 485.83789989989987u,0 486.8144399399399u,0 486.8154399399399u,1.5 487.79197997998u,1.5 487.79297997998u,0 488.7695200200201u,0 488.77052002002006u,1.5 489.7470600600601u,1.5 489.7480600600601u,0 495.6123003003003u,0 495.6133003003003u,1.5 497.56738038038037u,1.5 497.56838038038035u,0 499.5224604604605u,0 499.52346046046046u,1.5 500.5000005005005u,1.5 500.5010005005005u,0 503.4326206206207u,0 503.4336206206207u,1.5 504.41016066066067u,1.5 504.41116066066064u,0 507.34278078078074u,0 507.3437807807807u,1.5 508.3203208208209u,1.5 508.32132082082086u,0 509.2978608608609u,0 509.2988608608609u,1.5 510.2754009009009u,1.5 510.27640090090085u,0 518.0957212212213u,0 518.0967212212213u,1.5 519.0732612612613u,1.5 519.0742612612613u,0 521.0283413413413u,0 521.0293413413413u,1.5 522.0058813813813u,1.5 522.0068813813813u,0 525.9160415415415u,0 525.9170415415415u,1.5 526.8935815815815u,1.5 526.8945815815815u,0 528.8486616616617u,0 528.8496616616617u,1.5 530.8037417417418u,1.5 530.8047417417417u,0 531.7812817817818u,0 531.7822817817818u,1.5 533.7363618618618u,1.5 533.7373618618618u,0 534.7139019019019u,0 534.7149019019018u,1.5 540.5791421421421u,1.5 540.5801421421421u,0 542.5342222222223u,0 542.5352222222223u,1.5 545.4668423423423u,1.5 545.4678423423422u,0 546.4443823823824u,0 546.4453823823824u,1.5 547.4219224224224u,1.5 547.4229224224224u,0 548.3994624624625u,0 548.4004624624624u,1.5 549.3770025025025u,1.5 549.3780025025025u,0 550.3545425425425u,0 550.3555425425425u,1.5 551.3320825825826u,1.5 551.3330825825826u,0 553.2871626626627u,0 553.2881626626627u,1.5 554.2647027027027u,1.5 554.2657027027027u,0 560.1299429429429u,0 560.1309429429429u,1.5 561.107482982983u,1.5 561.108482982983u,0 563.0625630630631u,0 563.063563063063u,1.5 564.0401031031031u,1.5 564.0411031031031u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 569.9053433433434u,0 569.9063433433433u,1.5 575.7705835835836u,1.5 575.7715835835836u,0 576.7481236236237u,0 576.7491236236236u,1.5 577.7256636636637u,1.5 577.7266636636637u,0 584.5684439439439u,0 584.5694439439438u,1.5 585.545983983984u,1.5 585.546983983984u,0 587.501064064064u,0 587.502064064064u,1.5 589.4561441441441u,1.5 589.4571441441441u,0 590.4336841841842u,0 590.4346841841842u,1.5 592.3887642642643u,1.5 592.3897642642643u,0 594.3438443443445u,0 594.3448443443444u,1.5 595.3213843843844u,1.5 595.3223843843843u,0 598.2540045045045u,0 598.2550045045044u,1.5 599.2315445445446u,1.5 599.2325445445446u,0 600.2090845845846u,0 600.2100845845846u,1.5 601.1866246246246u,1.5 601.1876246246246u,0 602.1641646646647u,0 602.1651646646646u,1.5 603.1417047047047u,1.5 603.1427047047047u,0 605.0967847847849u,0 605.0977847847848u,1.5 606.0743248248249u,1.5 606.0753248248249u,0 607.0518648648649u,0 607.0528648648649u,1.5 613.8946451451452u,1.5 613.8956451451452u,0 615.8497252252253u,0 615.8507252252252u,1.5 616.8272652652653u,1.5 616.8282652652653u,0 620.7374254254254u,0 620.7384254254254u,1.5 621.7149654654654u,1.5 621.7159654654654u,0 623.6700455455456u,0 623.6710455455456u,1.5 628.5577457457458u,1.5 628.5587457457458u,0 637.355606106106u,0 637.356606106106u,1.5 643.2208463463464u,1.5 643.2218463463464u,0 645.1759264264264u,0 645.1769264264263u,1.5 646.1534664664664u,1.5 646.1544664664664u,0 649.0860865865866u,0 649.0870865865866u,1.5 653.9737867867868u,1.5 653.9747867867868u,0 654.9513268268269u,0 654.9523268268268u,1.5 656.9064069069069u,1.5 656.9074069069069u,0 660.816567067067u,0 660.817567067067u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 662.7716471471472u,0 662.7726471471472u,1.5 663.7491871871872u,1.5 663.7501871871872u,0 664.7267272272272u,0 664.7277272272272u,1.5 666.6818073073074u,1.5 666.6828073073074u,0 667.6593473473474u,0 667.6603473473474u,1.5 670.5919674674674u,1.5 670.5929674674674u,0 672.5470475475475u,0 672.5480475475475u,1.5 674.5021276276276u,1.5 674.5031276276276u,0 675.4796676676676u,0 675.4806676676676u,1.5 678.4122877877878u,1.5 678.4132877877878u,0 679.3898278278278u,0 679.3908278278278u,1.5 680.3673678678679u,1.5 680.3683678678678u,0 682.3224479479479u,0 682.3234479479479u,1.5 683.299987987988u,1.5 683.3009879879879u,0 685.255068068068u,0 685.256068068068u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 692.0978483483484u,1.5 692.0988483483484u,0 696.0080085085085u,0 696.0090085085085u,1.5 696.9855485485485u,1.5 696.9865485485485u,0 697.9630885885886u,0 697.9640885885885u,1.5 703.8283288288288u,1.5 703.8293288288288u,0 707.7384889889889u,0 707.7394889889889u,1.5 708.716029029029u,1.5 708.7170290290289u,0 709.693569069069u,0 709.694569069069u,1.5 712.6261891891892u,1.5 712.6271891891892u,0 713.6037292292292u,0 713.6047292292292u,1.5 714.5812692692692u,1.5 714.5822692692692u,0 716.5363493493494u,0 716.5373493493494u,1.5 717.5138893893894u,1.5 717.5148893893894u,0 718.4914294294294u,0 718.4924294294294u,1.5 722.4015895895895u,1.5 722.4025895895895u,0 723.3791296296296u,0 723.3801296296296u,1.5 724.3566696696697u,1.5 724.3576696696697u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 729.24436986987u,0 729.2453698698699u,1.5 730.22190990991u,1.5 730.22290990991u,0 731.19944994995u,0 731.20044994995u,1.5 733.15453003003u,1.5 733.1555300300299u,0 734.1320700700701u,0 734.1330700700701u,1.5 735.1096101101101u,1.5 735.1106101101101u,0 736.0871501501501u,0 736.0881501501501u,1.5 737.0646901901902u,1.5 737.0656901901901u,0 739.0197702702703u,0 739.0207702702703u,1.5 740.9748503503504u,1.5 740.9758503503504u,0 742.9299304304304u,0 742.9309304304304u,1.5 744.8850105105105u,1.5 744.8860105105105u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 755.637950950951u,1.5 755.638950950951u,0 756.615490990991u,0 756.616490990991u,1.5 757.593031031031u,1.5 757.594031031031u,0 764.4358113113113u,0 764.4368113113113u,1.5 765.4133513513514u,1.5 765.4143513513513u,0 766.3908913913914u,0 766.3918913913914u,1.5 767.3684314314314u,1.5 767.3694314314314u,0 770.3010515515515u,0 770.3020515515515u,1.5 771.2785915915915u,1.5 771.2795915915915u,0 772.2561316316315u,0 772.2571316316315u,1.5 775.1887517517517u,1.5 775.1897517517517u,0 776.1662917917918u,0 776.1672917917917u,1.5 777.1438318318318u,1.5 777.1448318318318u,0 781.053991991992u,0 781.054991991992u,1.5 782.031532032032u,1.5 782.032532032032u,0 783.0090720720721u,0 783.010072072072u,1.5 784.9641521521521u,1.5 784.9651521521521u,0 785.9416921921921u,0 785.9426921921921u,1.5 787.8967722722723u,1.5 787.8977722722723u,0 790.8293923923924u,0 790.8303923923924u,1.5 792.7844724724725u,1.5 792.7854724724725u,0 793.7620125125126u,0 793.7630125125125u,1.5 796.6946326326326u,1.5 796.6956326326326u,0 797.6721726726727u,0 797.6731726726726u,1.5 799.6272527527527u,1.5 799.6282527527527u,0 803.5374129129129u,0 803.5384129129129u,1.5 806.4700330330331u,1.5 806.4710330330331u,0 807.4475730730732u,0 807.4485730730731u,1.5 808.4251131131131u,1.5 808.426113113113u,0 814.2903533533533u,0 814.2913533533533u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 817.2229734734735u,0 817.2239734734735u,1.5 821.1331336336336u,1.5 821.1341336336336u,0 824.0657537537537u,0 824.0667537537537u,1.5 832.8636141141141u,1.5 832.864614114114u,0 835.7962342342342u,0 835.7972342342342u,1.5 836.7737742742743u,1.5 836.7747742742743u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 842.6390145145145u,0 842.6400145145145u,1.5 843.6165545545546u,1.5 843.6175545545545u,0 846.5491746746746u,0 846.5501746746746u,1.5 847.5267147147147u,1.5 847.5277147147146u,0 848.5042547547547u,0 848.5052547547547u,1.5 849.4817947947948u,1.5 849.4827947947948u,0 851.4368748748749u,0 851.4378748748749u,1.5 852.4144149149149u,1.5 852.4154149149149u,0 853.3919549549549u,0 853.3929549549549u,1.5 854.3694949949951u,1.5 854.370494994995u,0 859.2571951951952u,0 859.2581951951952u,1.5 860.2347352352352u,1.5 860.2357352352352u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 868.0550555555556u,1.5 868.0560555555555u,0 870.0101356356357u,0 870.0111356356357u,1.5 870.9876756756756u,1.5 870.9886756756756u,0 878.8079959959961u,0 878.808995995996u,1.5 882.7181561561562u,1.5 882.7191561561561u,0 883.6956961961962u,0 883.6966961961962u,1.5 886.6283163163163u,1.5 886.6293163163162u,0 894.4486366366367u,0 894.4496366366367u,1.5 896.4037167167166u,1.5 896.4047167167166u,0 897.3812567567567u,0 897.3822567567566u,1.5 902.2689569569569u,1.5 902.2699569569569u,0 904.2240370370371u,0 904.225037037037u,1.5 905.2015770770771u,1.5 905.2025770770771u,0 907.1566571571572u,0 907.1576571571571u,1.5 909.1117372372372u,1.5 909.1127372372372u,0 911.0668173173173u,0 911.0678173173172u,1.5 912.0443573573574u,1.5 912.0453573573574u,0 913.0218973973974u,0 913.0228973973974u,1.5 913.9994374374375u,1.5 914.0004374374374u,0 915.9545175175175u,0 915.9555175175175u,1.5 916.9320575575576u,1.5 916.9330575575576u,0 917.9095975975977u,0 917.9105975975976u,1.5 919.8646776776777u,1.5 919.8656776776777u,0 921.8197577577578u,0 921.8207577577577u,1.5 923.7748378378378u,1.5 923.7758378378378u,0 924.7523778778778u,0 924.7533778778778u,1.5 925.7299179179179u,1.5 925.7309179179178u,0 927.684997997998u,0 927.685997997998u,1.5 928.6625380380381u,1.5 928.663538038038u,0 932.5726981981983u,0 932.5736981981983u,1.5 933.5502382382382u,1.5 933.5512382382382u,0 935.5053183183182u,0 935.5063183183182u,1.5 938.4379384384384u,1.5 938.4389384384384u,0 939.4154784784785u,0 939.4164784784784u,1.5 947.2357987987988u,1.5 947.2367987987988u,0 948.2133388388388u,0 948.2143388388388u,1.5 949.1908788788788u,1.5 949.1918788788788u,0 950.1684189189189u,0 950.1694189189188u,1.5 951.145958958959u,1.5 951.146958958959u,0 957.0111991991993u,0 957.0121991991992u,1.5 957.9887392392392u,1.5 957.9897392392392u,0 959.9438193193192u,0 959.9448193193192u,1.5 960.9213593593594u,1.5 960.9223593593593u,0 964.8315195195195u,0 964.8325195195195u,1.5 966.7865995995996u,1.5 966.7875995995996u,0 967.7641396396397u,0 967.7651396396396u,1.5 968.7416796796797u,1.5 968.7426796796797u,0 970.6967597597597u,0 970.6977597597597u,1.5 972.6518398398398u,1.5 972.6528398398398u,0 973.6293798798798u,0 973.6303798798798u,1.5 974.60691991992u,1.5 974.6079199199199u,0 975.58445995996u,0 975.58545995996u,1.5 977.5395400400402u,1.5 977.5405400400401u,0 978.5170800800801u,0 978.51808008008u,1.5 981.4497002002003u,1.5 981.4507002002002u,0 984.3823203203203u,0 984.3833203203203u,1.5 986.3374004004004u,1.5 986.3384004004004u,0 987.3149404404405u,0 987.3159404404405u,1.5 989.2700205205206u,1.5 989.2710205205206u,0 992.2026406406408u,0 992.2036406406407u,1.5 993.1801806806807u,1.5 993.1811806806807u,0 995.1352607607607u,0 995.1362607607607u,1.5 999.045420920921u,1.5 999.0464209209209u,0 1000.0229609609609u,0 1000.0239609609608u,1.5 1001.9780410410411u,1.5 1001.9790410410411u,0 1002.955581081081u,0 1002.956581081081u,1.5 1003.9331211211212u,1.5 1003.9341211211212u,0 1005.8882012012012u,0 1005.8892012012012u,1.5 1006.8657412412414u,1.5 1006.8667412412414u,0 1007.8432812812813u,0 1007.8442812812813u,1.5 1013.7085215215216u,1.5 1013.7095215215215u,0 1014.6860615615615u,0 1014.6870615615614u,1.5 1016.6411416416418u,1.5 1016.6421416416417u,0 1017.6186816816817u,0 1017.6196816816816u,1.5 1021.5288418418419u,1.5 1021.5298418418419u,0 1022.5063818818818u,0 1022.5073818818818u,1.5 1026.416542042042u,1.5 1026.4175420420422u,0 1027.394082082082u,0 1027.3950820820821u,1.5 1028.371622122122u,1.5 1028.3726221221223u,0 1029.349162162162u,0 1029.3501621621622u,1.5 1030.3267022022021u,1.5 1030.3277022022023u,0 1031.3042422422423u,0 1031.3052422422425u,1.5 1032.2817822822822u,1.5 1032.2827822822824u,0 1033.2593223223223u,0 1033.2603223223225u,1.5 1034.2368623623622u,1.5 1034.2378623623624u,0 1041.0796426426425u,0 1041.0806426426427u,1.5 1042.0571826826824u,1.5 1042.0581826826826u,0 1045.9673428428428u,0 1045.968342842843u,1.5 1046.9448828828827u,1.5 1046.9458828828829u,0 1047.9224229229228u,0 1047.923422922923u,1.5 1048.8999629629627u,1.5 1048.900962962963u,0 1049.8775030030029u,0 1049.878503003003u,1.5 1050.855043043043u,1.5 1050.8560430430432u,0 1051.832583083083u,0 1051.833583083083u,1.5 1052.810123123123u,1.5 1052.8111231231233u,0 1053.787663163163u,0 1053.7886631631632u,1.5 1054.765203203203u,1.5 1054.7662032032033u,0 1055.7427432432432u,0 1055.7437432432434u,1.5 1057.6978233233233u,1.5 1057.6988233233235u,0 1058.6753633633632u,0 1058.6763633633634u,1.5 1061.6079834834834u,1.5 1061.6089834834836u,0 1062.5855235235235u,0 1062.5865235235237u,1.5 1065.5181436436435u,1.5 1065.5191436436437u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1070.4058438438437u,0 1070.406843843844u,1.5 1071.3833838838837u,1.5 1071.3843838838839u,0 1077.248624124124u,0 1077.2496241241242u,1.5 1079.203704204204u,1.5 1079.2047042042043u,0 1080.1812442442442u,0 1080.1822442442444u,1.5 1081.1587842842841u,1.5 1081.1597842842843u,0 1082.1363243243243u,0 1082.1373243243245u,1.5 1086.0464844844844u,1.5 1086.0474844844846u,0 1087.0240245245245u,0 1087.0250245245247u,1.5 1093.8668048048046u,1.5 1093.8678048048048u,0 1096.7994249249248u,0 1096.800424924925u,1.5 1102.6646651651652u,1.5 1102.6656651651654u,0 1103.642205205205u,0 1103.6432052052053u,1.5 1104.6197452452452u,1.5 1104.6207452452454u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1107.5523653653654u,1.5 1107.5533653653656u,0 1108.5299054054053u,0 1108.5309054054055u,1.5 1109.5074454454455u,1.5 1109.5084454454457u,0 1113.4176056056056u,0 1113.4186056056058u,1.5 1115.3726856856854u,1.5 1115.3736856856856u,0 1116.3502257257255u,0 1116.3512257257257u,1.5 1119.2828458458457u,1.5 1119.283845845846u,0 1121.2379259259258u,0 1121.238925925926u,1.5 1122.215465965966u,1.5 1122.216465965966u,0 1124.170546046046u,0 1124.1715460460462u,1.5 1125.1480860860859u,1.5 1125.149086086086u,0 1126.125626126126u,0 1126.1266261261262u,1.5 1127.1031661661661u,1.5 1127.1041661661664u,0 1130.035786286286u,0 1130.0367862862863u,1.5 1131.0133263263263u,1.5 1131.0143263263265u,0 1131.9908663663664u,0 1131.9918663663666u,1.5 1134.9234864864864u,1.5 1134.9244864864866u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1142.7438068068066u,0 1142.7448068068068u,1.5 1143.7213468468467u,1.5 1143.722346846847u,0 1144.6988868868866u,0 1144.6998868868868u,1.5 1148.609047047047u,1.5 1148.6100470470471u,0 1150.564127127127u,0 1150.5651271271272u,1.5 1156.4293673673674u,1.5 1156.4303673673676u,0 1158.3844474474474u,0 1158.3854474474476u,1.5 1161.3170675675676u,1.5 1161.3180675675678u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1165.2272277277275u,1.5 1165.2282277277277u,0 1166.2047677677676u,0 1166.2057677677678u,1.5 1167.1823078078075u,1.5 1167.1833078078078u,0 1170.1149279279277u,0 1170.115927927928u,1.5 1172.0700080080078u,1.5 1172.071008008008u,0 1173.047548048048u,0 1173.0485480480481u,1.5 1175.002628128128u,1.5 1175.0036281281282u,0 1176.957708208208u,0 1176.9587082082082u,1.5 1178.912788288288u,1.5 1178.9137882882883u,0 1179.8903283283282u,0 1179.8913283283284u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1190.6432687687686u,0 1190.6442687687688u,1.5 1191.6208088088085u,1.5 1191.6218088088087u,0 1192.5983488488487u,0 1192.5993488488489u,1.5 1197.486049049049u,1.5 1197.4870490490491u,0 1199.441129129129u,0 1199.4421291291292u,1.5 1200.418669169169u,1.5 1200.4196691691693u,0 1201.396209209209u,0 1201.3972092092092u,1.5 1202.3737492492492u,1.5 1202.3747492492494u,0 1203.3512892892893u,0 1203.3522892892895u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1208.2389894894895u,0 1208.2399894894897u,1.5 1210.1940695695696u,1.5 1210.1950695695698u,0 1213.1266896896898u,0 1213.12768968969u,1.5 1214.1042297297297u,1.5 1214.10522972973u,0 1215.0817697697696u,0 1215.0827697697698u,1.5 1217.0368498498497u,1.5 1217.0378498498499u,0 1218.0143898898898u,0 1218.01538988989u,1.5 1218.9919299299297u,1.5 1218.99292992993u,0 1219.9694699699699u,0 1219.97046996997u,1.5 1220.9470100100098u,1.5 1220.94801001001u,0 1223.87963013013u,0 1223.8806301301302u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1232.6774904904905u,1.5 1232.6784904904907u,0 1234.6325705705706u,0 1234.6335705705708u,1.5 1241.4753508508506u,1.5 1241.4763508508508u,0 1242.4528908908908u,0 1242.453890890891u,1.5 1243.4304309309307u,1.5 1243.431430930931u,0 1244.4079709709708u,0 1244.408970970971u,1.5 1245.3855110110107u,1.5 1245.386511011011u,0 1246.363051051051u,0 1246.364051051051u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1260.0486116116115u,1.5 1260.0496116116117u,0 1261.0261516516516u,0 1261.0271516516518u,1.5 1262.0036916916918u,1.5 1262.004691691692u,0 1265.9138518518516u,0 1265.9148518518518u,1.5 1266.8913918918918u,1.5 1266.892391891892u,0 1267.8689319319317u,0 1267.869931931932u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1271.779092092092u,0 1271.7800920920922u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1276.6667922922923u,0 1276.6677922922925u,1.5 1278.6218723723723u,1.5 1278.6228723723725u,0 1279.5994124124122u,0 1279.6004124124124u,1.5 1280.5769524524524u,1.5 1280.5779524524526u,0 1287.4197327327327u,0 1287.4207327327329u,1.5 1288.3972727727728u,1.5 1288.398272772773u,0 1289.3748128128127u,0 1289.375812812813u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1291.3298928928928u,0 1291.330892892893u,1.5 1292.3074329329327u,1.5 1292.3084329329329u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1295.2400530530529u,1.5 1295.241053053053u,0 1298.172673173173u,0 1298.1736731731733u,1.5 1303.0603733733733u,1.5 1303.0613733733735u,0 1305.0154534534533u,0 1305.0164534534536u,1.5 1305.9929934934935u,1.5 1305.9939934934937u,0 1306.9705335335334u,0 1306.9715335335336u,1.5 1307.9480735735735u,1.5 1307.9490735735737u,0 1308.9256136136135u,0 1308.9266136136137u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1315.7683938938937u,0 1315.769393893894u,1.5 1316.7459339339337u,1.5 1316.7469339339339u,0 1318.701014014014u,0 1318.7020140140141u,1.5 1319.6785540540538u,1.5 1319.679554054054u,0 1320.656094094094u,0 1320.6570940940942u,1.5 1327.4988743743743u,1.5 1327.4998743743745u,0 1329.4539544544543u,0 1329.4549544544545u,1.5 1332.3865745745745u,1.5 1332.3875745745747u,0 1333.3641146146147u,0 1333.3651146146149u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1343.139515015015u,1.5 1343.1405150150151u,0 1344.1170550550548u,0 1344.118055055055u,1.5 1345.094595095095u,1.5 1345.0955950950952u,0 1346.0721351351349u,0 1346.073135135135u,1.5 1347.049675175175u,1.5 1347.0506751751752u,0 1349.004755255255u,0 1349.0057552552553u,1.5 1350.9598353353351u,1.5 1350.9608353353353u,0 1352.9149154154154u,0 1352.9159154154156u,1.5 1353.8924554554553u,1.5 1353.8934554554555u,0 1356.8250755755755u,0 1356.8260755755757u,1.5 1358.7801556556556u,1.5 1358.7811556556558u,0 1359.7576956956957u,0 1359.758695695696u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1367.578016016016u,0 1367.579016016016u,1.5 1368.5555560560558u,1.5 1368.556556056056u,0 1369.533096096096u,0 1369.5340960960962u,1.5 1370.5106361361359u,1.5 1370.511636136136u,0 1371.488176176176u,0 1371.4891761761762u,1.5 1373.443256256256u,1.5 1373.4442562562563u,0 1374.4207962962962u,0 1374.4217962962964u,1.5 1376.3758763763763u,1.5 1376.3768763763765u,0 1377.3534164164164u,0 1377.3544164164166u,1.5 1378.3309564564563u,1.5 1378.3319564564565u,0 1379.3084964964964u,0 1379.3094964964966u,1.5 1380.2860365365364u,1.5 1380.2870365365366u,0 1383.2186566566565u,0 1383.2196566566568u,1.5 1385.1737367367366u,1.5 1385.1747367367368u,0 1386.1512767767767u,0 1386.152276776777u,1.5 1387.1288168168169u,1.5 1387.129816816817u,0 1388.1063568568568u,0 1388.107356856857u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1399.836837337337u,0 1399.8378373373373u,1.5 1403.7469974974974u,1.5 1403.7479974974976u,0 1404.7245375375373u,0 1404.7255375375375u,1.5 1406.6796176176176u,1.5 1406.6806176176178u,0 1407.6571576576575u,0 1407.6581576576577u,1.5 1408.6346976976977u,1.5 1408.6356976976979u,0 1409.6122377377376u,0 1409.6132377377378u,1.5 1411.5673178178179u,1.5 1411.568317817818u,0 1414.4999379379378u,0 1414.500937937938u,1.5 1415.4774779779777u,1.5 1415.478477977978u,0 1418.410098098098u,0 1418.4110980980981u,1.5 1419.3876381381378u,1.5 1419.388638138138u,0 1420.365178178178u,0 1420.3661781781782u,1.5 1421.3427182182181u,1.5 1421.3437182182183u,0 1422.320258258258u,0 1422.3212582582582u,1.5 1423.2977982982982u,1.5 1423.2987982982984u,0 1425.2528783783782u,0 1425.2538783783784u,1.5 1426.2304184184184u,1.5 1426.2314184184186u,0 1427.2079584584583u,0 1427.2089584584585u,1.5 1430.1405785785785u,1.5 1430.1415785785787u,0 1432.0956586586585u,0 1432.0966586586587u,1.5 1433.0731986986987u,1.5 1433.0741986986989u,0 1434.0507387387386u,0 1434.0517387387388u,1.5 1436.0058188188189u,1.5 1436.006818818819u,0 1438.938438938939u,0 1438.9394389389392u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1440.8935190190189u,0 1440.894519019019u,1.5 1441.8710590590588u,1.5 1441.872059059059u,0 1444.803679179179u,0 1444.8046791791792u,1.5 1445.781219219219u,1.5 1445.7822192192193u,0 1446.758759259259u,0 1446.7597592592592u,1.5 1447.7362992992992u,1.5 1447.7372992992994u,0 1449.6913793793792u,0 1449.6923793793794u,1.5 1450.6689194194194u,1.5 1450.6699194194196u,0 1451.6464594594593u,0 1451.6474594594595u,1.5 1453.6015395395395u,1.5 1453.6025395395397u,0 1454.5790795795795u,0 1454.5800795795797u,1.5 1464.35447997998u,1.5 1464.3554799799801u,0 1465.3320200200199u,0 1465.33302002002u,1.5 1467.2871001001u,1.5 1467.2881001001u,0 1468.26464014014u,0 1468.2656401401402u,1.5 1470.21972022022u,1.5 1470.2207202202203u,0 1471.19726026026u,0 1471.1982602602602u,1.5 1473.1523403403403u,1.5 1473.1533403403405u,0 1474.1298803803802u,0 1474.1308803803804u,1.5 1476.0849604604603u,1.5 1476.0859604604605u,0 1477.0625005005004u,0 1477.0635005005006u,1.5 1478.0400405405405u,1.5 1478.0410405405407u,0 1480.9726606606605u,0 1480.9736606606607u,1.5 1481.9502007007006u,1.5 1481.9512007007008u,0 1482.9277407407408u,0 1482.928740740741u,1.5 1483.9052807807807u,1.5 1483.906280780781u,0 1489.7705210210208u,0 1489.771521021021u,1.5 1490.7480610610608u,1.5 1490.749061061061u,0 1494.658221221221u,0 1494.6592212212213u,1.5 1495.635761261261u,1.5 1495.6367612612612u,0 1510.2988618618617u,0 1510.299861861862u,1.5 1511.2764019019019u,1.5 1511.277401901902u,0 1513.231481981982u,0 1513.2324819819821u,1.5 1514.209022022022u,1.5 1514.2100220220223u,0 1518.119182182182u,0 1518.1201821821821u,1.5 1519.096722222222u,1.5 1519.0977222222223u,0 1520.074262262262u,0 1520.0752622622622u,1.5 1521.0518023023021u,1.5 1521.0528023023023u,0 1522.0293423423423u,0 1522.0303423423425u,1.5 1523.0068823823822u,1.5 1523.0078823823824u,0 1524.9619624624622u,0 1524.9629624624624u,1.5 1525.9395025025024u,1.5 1525.9405025025026u,0 1526.9170425425425u,0 1526.9180425425427u,1.5 1527.8945825825824u,1.5 1527.8955825825826u,0 1530.8272027027026u,0 1530.8282027027028u,1.5 1531.8047427427427u,1.5 1531.805742742743u,0 1532.7822827827827u,0 1532.7832827827829u,1.5 1542.557683183183u,1.5 1542.5586831831831u,0 1543.535223223223u,0 1543.5362232232233u,1.5 1545.490303303303u,1.5 1545.4913033033033u,0 1546.4678433433432u,0 1546.4688433433435u,1.5 1548.4229234234233u,1.5 1548.4239234234235u,0 1549.4004634634632u,0 1549.4014634634634u,1.5 1550.3780035035034u,1.5 1550.3790035035036u,0 1551.3555435435435u,0 1551.3565435435437u,1.5 1552.3330835835834u,1.5 1552.3340835835836u,0 1553.3106236236235u,0 1553.3116236236237u,1.5 1554.2881636636635u,1.5 1554.2891636636637u,0 1562.108483983984u,0 1562.109483983984u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1565.041104104104u,0 1565.0421041041043u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1567.973724224224u,0 1567.9747242242242u,1.5 1575.7940445445445u,1.5 1575.7950445445447u,0 1576.7715845845844u,0 1576.7725845845846u,1.5 1582.6368248248248u,1.5 1582.637824824825u,0 1583.614364864865u,0 1583.6153648648651u,1.5 1585.569444944945u,1.5 1585.5704449449452u,0 1586.5469849849849u,0 1586.547984984985u,1.5 1587.524525025025u,1.5 1587.5255250250252u,0 1589.479605105105u,0 1589.4806051051053u,1.5 1596.3223853853851u,1.5 1596.3233853853853u,0 1597.2999254254253u,0 1597.3009254254255u,1.5 1598.2774654654654u,1.5 1598.2784654654656u,0 1601.2100855855854u,0 1601.2110855855856u,1.5 1603.1651656656657u,1.5 1603.1661656656659u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1607.0753258258258u,0 1607.076325825826u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1613.918106106106u,1.5 1613.9191061061063u,0 1618.805806306306u,0 1618.8068063063063u,1.5 1619.7833463463462u,1.5 1619.7843463463464u,0 1621.7384264264263u,0 1621.7394264264265u,1.5 1628.5812067067066u,1.5 1628.5822067067068u,0 1629.5587467467467u,0 1629.559746746747u,1.5 1630.5362867867866u,1.5 1630.5372867867868u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1641.289227227227u,1.5 1641.2902272272272u,0 1642.2667672672671u,0 1642.2677672672673u,1.5 1643.244307307307u,1.5 1643.2453073073073u,0 1644.2218473473472u,0 1644.2228473473474u,1.5 1645.199387387387u,1.5 1645.2003873873873u,0 1650.0870875875873u,0 1650.0880875875876u,1.5 1651.0646276276275u,1.5 1651.0656276276277u,0 1652.0421676676676u,0 1652.0431676676678u,1.5 1654.9747877877876u,1.5 1654.9757877877878u,0 1656.9298678678679u,0 1656.930867867868u,1.5 1657.9074079079078u,1.5 1657.908407907908u,0 1662.795108108108u,0 1662.7961081081082u,1.5 1665.727728228228u,1.5 1665.7287282282282u,0 1666.7052682682681u,0 1666.7062682682683u,1.5 1668.6603483483482u,1.5 1668.6613483483484u,0 1674.5255885885883u,0 1674.5265885885885u,1.5 1675.5031286286285u,1.5 1675.5041286286287u,0 1677.4582087087085u,0 1677.4592087087087u,1.5 1678.4357487487487u,1.5 1678.4367487487489u,0 1679.4132887887886u,0 1679.4142887887888u,1.5 1680.3908288288287u,1.5 1680.391828828829u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1689.1886891891893u,1.5 1689.1896891891895u,0 1691.1437692692691u,0 1691.1447692692693u,1.5 1693.0988493493492u,1.5 1693.0998493493494u,0 1695.0539294294292u,0 1695.0549294294294u,1.5 1696.0314694694694u,1.5 1696.0324694694696u,0 1698.9640895895895u,0 1698.9650895895898u,1.5 1701.8967097097095u,1.5 1701.8977097097097u,0 1702.8742497497497u,0 1702.8752497497499u,1.5 1705.8068698698698u,1.5 1705.80786986987u,0 1707.76194994995u,0 1707.76294994995u,1.5 1712.6496501501501u,1.5 1712.6506501501503u,0 1713.6271901901903u,0 1713.6281901901905u,1.5 1714.6047302302302u,1.5 1714.6057302302304u,0 1719.4924304304302u,0 1719.4934304304304u,1.5 1720.4699704704703u,1.5 1720.4709704704705u,0 1721.4475105105103u,0 1721.4485105105105u,1.5 1723.4025905905905u,1.5 1723.4035905905907u,0 1727.3127507507506u,0 1727.3137507507508u,1.5 1729.2678308308307u,1.5 1729.268830830831u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1735.133071071071u,1.5 1735.1340710710713u,0 1737.0881511511511u,0 1737.0891511511513u,1.5 1738.0656911911913u,1.5 1738.0666911911915u,0 1740.998311311311u,0 1740.9993113113112u,1.5 1741.9758513513511u,1.5 1741.9768513513513u,0 1742.9533913913913u,0 1742.9543913913915u,1.5 1745.8860115115112u,1.5 1745.8870115115114u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1754.6838718718718u,0 1754.684871871872u,1.5 1755.6614119119117u,1.5 1755.662411911912u,0 1758.594032032032u,0 1758.5950320320321u,1.5 1759.571572072072u,1.5 1759.5725720720723u,0 1761.526652152152u,0 1761.5276521521523u,1.5 1764.4592722722723u,1.5 1764.4602722722725u,0 1766.4143523523521u,0 1766.4153523523523u,1.5 1768.3694324324322u,1.5 1768.3704324324324u,0 1771.3020525525524u,0 1771.3030525525526u,1.5 1774.2346726726726u,1.5 1774.2356726726728u,0 1775.2122127127125u,0 1775.2132127127127u,1.5 1777.1672927927928u,1.5 1777.168292792793u,0 1779.1223728728728u,0 1779.123372872873u,1.5 1780.0999129129127u,1.5 1780.100912912913u,0 1781.0774529529529u,0 1781.078452952953u,1.5 1784.010073073073u,1.5 1784.0110730730732u,0 1784.987613113113u,0 1784.9886131131132u,1.5 1788.8977732732733u,1.5 1788.8987732732735u,0 1790.852853353353u,0 1790.8538533533533u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1794.7630135135132u,1.5 1794.7640135135134u,0 1796.7180935935935u,0 1796.7190935935937u,1.5 1798.6731736736735u,1.5 1798.6741736736737u,0 1802.5833338338336u,0 1802.5843338338339u,1.5 1803.5608738738738u,1.5 1803.561873873874u,0 1804.5384139139137u,0 1804.539413913914u,1.5 1807.471034034034u,1.5 1807.472034034034u,0 1808.448574074074u,0 1808.4495740740742u,1.5 1809.426114114114u,1.5 1809.4271141141141u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1820.1790545545543u,1.5 1820.1800545545545u,0 1821.1565945945945u,0 1821.1575945945947u,1.5 1822.1341346346344u,1.5 1822.1351346346346u,0 1823.1116746746745u,0 1823.1126746746747u,1.5 1824.0892147147147u,1.5 1824.0902147147149u,0 1826.0442947947947u,0 1826.045294794795u,1.5 1832.887075075075u,1.5 1832.8880750750752u,0 1834.842155155155u,0 1834.8431551551553u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1839.7298553553553u,0 1839.7308553553555u,1.5 1843.6400155155154u,1.5 1843.6410155155156u,0 1845.5950955955955u,0 1845.5960955955957u,1.5 1846.5726356356354u,1.5 1846.5736356356356u,0 1851.4603358358356u,0 1851.4613358358358u,1.5 1854.3929559559558u,1.5 1854.393955955956u,0 1857.325576076076u,0 1857.3265760760762u,1.5 1858.3031161161161u,1.5 1858.3041161161163u,0 1863.1908163163164u,0 1863.1918163163166u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1866.1234364364361u,0 1866.1244364364363u,1.5 1871.0111366366364u,1.5 1871.0121366366366u,0 1871.9886766766765u,0 1871.9896766766767u,1.5 1872.9662167167166u,1.5 1872.9672167167168u,0 1876.8763768768767u,0 1876.877376876877u,1.5 1877.853916916917u,1.5 1877.854916916917u,0 1878.8314569569568u,0 1878.832456956957u,1.5 1883.719157157157u,1.5 1883.7201571571572u,0 1884.6966971971972u,0 1884.6976971971974u,1.5 1885.674237237237u,1.5 1885.6752372372373u,0 1887.6293173173174u,0 1887.6303173173176u,1.5 1888.6068573573573u,1.5 1888.6078573573575u,0 1889.5843973973974u,0 1889.5853973973976u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1900.3373378378376u,0 1900.3383378378378u,1.5 1903.2699579579578u,1.5 1903.270957957958u,0 1905.2250380380378u,0 1905.226038038038u,1.5 1906.202578078078u,1.5 1906.2035780780782u,0 1908.157658158158u,0 1908.1586581581582u,1.5 1909.1351981981982u,1.5 1909.1361981981984u,0 1911.0902782782782u,0 1911.0912782782784u,1.5 1915.0004384384383u,1.5 1915.0014384384385u,0 1916.9555185185184u,0 1916.9565185185186u,1.5 1919.8881386386383u,1.5 1919.8891386386385u,0 1920.8656786786785u,0 1920.8666786786787u,1.5 1922.8207587587585u,1.5 1922.8217587587587u,0 1924.7758388388386u,0 1924.7768388388388u,1.5 1925.7533788788787u,1.5 1925.754378878879u,0 1926.7309189189189u,0 1926.731918918919u,1.5 1927.7084589589588u,1.5 1927.709458958959u,0 1929.6635390390388u,0 1929.664539039039u,1.5 1930.641079079079u,1.5 1930.6420790790792u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1940.4164794794794u,1.5 1940.4174794794797u,0 1942.3715595595593u,0 1942.3725595595595u,1.5 1943.3490995995994u,1.5 1943.3500995995996u,0 1946.2817197197196u,0 1946.2827197197198u,1.5 1948.2367997997997u,1.5 1948.2377997997999u,0 1949.2143398398398u,0 1949.21533983984u,1.5 1950.1918798798797u,1.5 1950.19287987988u,0 1951.1694199199198u,0 1951.17041991992u,1.5 1953.1245u,1.5 1953.1255u,0 1956.0571201201199u,0 1956.05812012012u,1.5 1957.03466016016u,1.5 1957.0356601601602u,0 1958.9897402402403u,0 1958.9907402402405u,1.5 1961.9223603603602u,1.5 1961.9233603603604u,0 1964.8549804804804u,0 1964.8559804804806u,1.5 1965.8325205205203u,1.5 1965.8335205205206u,0 1967.7876006006004u,0 1967.7886006006006u,1.5 1968.7651406406405u,1.5 1968.7661406406407u,0 1970.7202207207204u,0 1970.7212207207206u,1.5 1971.6977607607605u,1.5 1971.6987607607607u,0 1974.630380880881u,0 1974.6313808808811u,1.5 1976.5854609609607u,1.5 1976.586460960961u,0 1977.5630010010009u,0 1977.564001001001u,1.5 1980.4956211211208u,1.5 1980.496621121121u,0 1981.473161161161u,0 1981.4741611611612u,1.5 1983.4282412412413u,1.5 1983.4292412412415u,0 1984.4057812812814u,0 1984.4067812812816u,1.5 1986.3608613613612u,1.5 1986.3618613613614u,0 1991.2485615615612u,0 1991.2495615615614u,1.5 1992.2261016016014u,1.5 1992.2271016016016u,0 1993.2036416416415u,0 1993.2046416416417u,1.5 1995.1587217217213u,1.5 1995.1597217217216u,0 1997.1138018018016u,0 1997.1148018018018u,1.5 1998.0913418418418u,1.5 1998.092341841842u,0 1999.068881881882u,0 1999.069881881882u,1.5 2005.911662162162u,1.5 2005.9126621621622u,0 2006.8892022022021u,0 2006.8902022022023u,1.5 2007.8667422422423u,1.5 2007.8677422422425u,0 2009.821822322322u,0 2009.8228223223223u,1.5 2014.7095225225223u,1.5 2014.7105225225225u,0 2015.6870625625625u,0 2015.6880625625627u,1.5 2021.5523028028026u,1.5 2021.5533028028028u,0 2022.5298428428428u,0 2022.530842842843u,1.5 2023.507382882883u,1.5 2023.508382882883u,0 2024.4849229229226u,0 2024.4859229229228u,1.5 2025.4624629629627u,1.5 2025.463462962963u,0 2026.4400030030029u,0 2026.441003003003u,1.5 2027.417543043043u,1.5 2027.4185430430432u,0 2028.3950830830831u,0 2028.3960830830833u,1.5 2029.3726231231228u,1.5 2029.373623123123u,0 2032.3052432432432u,0 2032.3062432432434u,1.5 2033.2827832832834u,1.5 2033.2837832832836u,0 2036.2154034034033u,0 2036.2164034034035u,1.5 2037.1929434434435u,1.5 2037.1939434434437u,0 2040.1255635635634u,0 2040.1265635635636u,1.5 2042.0806436436435u,1.5 2042.0816436436437u,0 2043.0581836836836u,0 2043.0591836836838u,1.5 2044.0357237237233u,1.5 2044.0367237237235u,0 2046.9683438438437u,0 2046.969343843844u,1.5 2047.9458838838839u,1.5 2047.946883883884u,0 2048.9234239239236u,0 2048.9244239239238u,1.5 2049.900963963964u,1.5 2049.901963963964u,0 2051.856044044044u,0 2051.8570440440444u,1.5 2054.788664164164u,1.5 2054.789664164164u,0 2055.766204204204u,0 2055.767204204204u,1.5 2058.698824324324u,1.5 2058.6998243243243u,0 2060.6539044044043u,0 2060.6549044044045u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2067.4966846846846u,1.5 2067.497684684685u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2070.429304804805u,1.5 2070.430304804805u,0 2074.339464964965u,0 2074.340464964965u,1.5 2075.317005005005u,1.5 2075.318005005005u,0 2077.272085085085u,0 2077.2730850850853u,1.5 2078.249625125125u,1.5 2078.250625125125u,0 2079.227165165165u,0 2079.228165165165u,1.5 2086.0699454454452u,1.5 2086.0709454454454u,0 2091.9351856856856u,0 2091.936185685686u,1.5 2092.9127257257255u,1.5 2092.9137257257257u,0 2095.8453458458457u,0 2095.846345845846u,1.5 2096.822885885886u,1.5 2096.8238858858863u,0 2097.8004259259255u,0 2097.8014259259257u,1.5 2102.688126126126u,1.5 2102.689126126126u,0 2104.643206206206u,0 2104.644206206206u,1.5 2105.620746246246u,1.5 2105.6217462462464u,0 2114.4186066066063u,0 2114.4196066066065u,1.5 2120.2838468468467u,1.5 2120.284846846847u,0 2121.261386886887u,0 2121.2623868868873u,1.5 2123.216466966967u,1.5 2123.217466966967u,0 2127.126627127127u,0 2127.127627127127u,1.5 2128.104167167167u,1.5 2128.105167167167u,0 2129.081707207207u,0 2129.082707207207u,1.5 2132.991867367367u,1.5 2132.992867367367u,0 2133.9694074074073u,0 2133.9704074074075u,1.5 2134.946947447447u,1.5 2134.9479474474474u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2137.8795675675674u,1.5 2137.8805675675676u,0 2138.8571076076073u,0 2138.8581076076075u,1.5 2140.8121876876876u,1.5 2140.813187687688u,0 2142.7672677677674u,0 2142.7682677677676u,1.5 2143.744807807808u,1.5 2143.745807807808u,0 2144.7223478478477u,0 2144.723347847848u,1.5 2145.699887887888u,1.5 2145.7008878878883u,0 2146.677427927928u,0 2146.678427927928u,1.5 2149.610048048048u,1.5 2149.6110480480484u,0 2154.497748248248u,0 2154.4987482482484u,1.5 2156.4528283283285u,1.5 2156.4538283283287u,0 2157.430368368368u,0 2157.431368368368u,1.5 2162.3180685685684u,1.5 2162.3190685685686u,0 2163.2956086086083u,0 2163.2966086086085u,1.5 2164.2731486486487u,1.5 2164.274148648649u,0 2167.2057687687684u,0 2167.2067687687686u,1.5 2169.1608488488487u,1.5 2169.161848848849u,0 2170.138388888889u,0 2170.1393888888892u,1.5 2174.048549049049u,1.5 2174.0495490490493u,0 2180.8913293293294u,0 2180.8923293293296u,1.5 2181.868869369369u,1.5 2181.869869369369u,0 2182.8464094094093u,0 2182.8474094094095u,1.5 2184.8014894894895u,1.5 2184.8024894894897u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2187.7341096096093u,1.5 2187.7351096096095u,0 2191.6442697697694u,0 2191.6452697697696u,1.5 2196.53196996997u,1.5 2196.53296996997u,0 2197.5095100100098u,0 2197.51051001001u,1.5 2198.48705005005u,1.5 2198.4880500500503u,0 2200.4421301301304u,0 2200.4431301301306u,1.5 2201.41967017017u,1.5 2201.42067017017u,0 2203.37475025025u,0 2203.3757502502503u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2211.1950705705704u,0 2211.1960705705706u,1.5 2212.1726106106103u,1.5 2212.1736106106105u,0 2215.105230730731u,0 2215.106230730731u,1.5 2219.992930930931u,1.5 2219.993930930931u,0 2220.970470970971u,0 2220.971470970971u,1.5 2221.9480110110107u,1.5 2221.949011011011u,0 2223.903091091091u,0 2223.9040910910912u,1.5 2227.813251251251u,1.5 2227.8142512512513u,0 2228.790791291291u,0 2228.7917912912912u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2230.745871371371u,0 2230.746871371371u,1.5 2232.700951451451u,1.5 2232.7019514514514u,0 2234.6560315315314u,0 2234.6570315315316u,1.5 2235.6335715715713u,1.5 2235.6345715715715u,0 2236.6111116116112u,0 2236.6121116116115u,1.5 2238.5661916916915u,1.5 2238.5671916916917u,0 2239.543731731732u,0 2239.544731731732u,1.5 2240.5212717717714u,1.5 2240.5222717717716u,0 2241.4988118118117u,0 2241.499811811812u,1.5 2242.4763518518516u,1.5 2242.477351851852u,0 2243.453891891892u,0 2243.454891891892u,1.5 2244.431431931932u,1.5 2244.432431931932u,0 2245.408971971972u,0 2245.409971971972u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2255.184372372372u,1.5 2255.185372372372u,0 2256.161912412412u,0 2256.1629124124124u,1.5 2260.0720725725723u,1.5 2260.0730725725725u,0 2264.9597727727723u,0 2264.9607727727725u,1.5 2265.9373128128127u,1.5 2265.938312812813u,0 2266.9148528528526u,0 2266.915852852853u,1.5 2267.892392892893u,1.5 2267.893392892893u,0 2269.847472972973u,0 2269.848472972973u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2276.690253253253u,0 2276.6912532532533u,1.5 2277.6677932932935u,1.5 2277.6687932932937u,0 2278.6453333333334u,0 2278.6463333333336u,1.5 2280.600413413413u,1.5 2280.6014134134134u,0 2281.577953453453u,0 2281.5789534534533u,1.5 2282.5554934934935u,1.5 2282.5564934934937u,0 2284.5105735735733u,0 2284.5115735735735u,1.5 2285.488113613613u,1.5 2285.4891136136134u,0 2287.4431936936935u,0 2287.4441936936937u,1.5 2288.420733733734u,1.5 2288.421733733734u,0 2289.3982737737733u,0 2289.3992737737735u,1.5 2290.3758138138137u,1.5 2290.376813813814u,0 2292.330893893894u,0 2292.331893893894u,1.5 2293.308433933934u,1.5 2293.309433933934u,0 2299.173674174174u,0 2299.174674174174u,1.5 2304.0613743743743u,1.5 2304.0623743743745u,0 2307.9715345345344u,0 2307.9725345345346u,1.5 2308.9490745745743u,1.5 2308.9500745745745u,0 2309.926614614614u,0 2309.9276146146144u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2314.8143148148147u,0 2314.815314814815u,1.5 2319.7020150150147u,1.5 2319.703015015015u,0 2320.679555055055u,0 2320.6805550550553u,1.5 2324.589715215215u,1.5 2324.5907152152154u,0 2325.567255255255u,0 2325.5682552552553u,1.5 2327.5223353353354u,1.5 2327.5233353353356u,0 2332.4100355355354u,0 2332.4110355355356u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2340.2303558558556u,0 2340.231355855856u,1.5 2341.207895895896u,1.5 2341.208895895896u,0 2342.185435935936u,0 2342.186435935936u,1.5 2343.1629759759758u,1.5 2343.163975975976u,0 2344.1405160160157u,0 2344.141516016016u,1.5 2349.028216216216u,1.5 2349.0292162162164u,0 2350.005756256256u,0 2350.0067562562563u,1.5 2350.9832962962964u,1.5 2350.9842962962966u,0 2354.893456456456u,0 2354.8944564564563u,1.5 2355.8709964964964u,1.5 2355.8719964964966u,0 2356.8485365365364u,0 2356.8495365365366u,1.5 2358.803616616616u,1.5 2358.8046166166164u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2366.623936936937u,1.5 2366.624936936937u,0 2367.6014769769768u,0 2367.602476976977u,1.5 2369.556557057057u,1.5 2369.5575570570572u,0 2371.5116371371373u,0 2371.5126371371375u,1.5 2376.3993373373373u,1.5 2376.4003373373375u,0 2377.3768773773777u,0 2377.377877377378u,1.5 2380.3094974974974u,1.5 2380.3104974974976u,0 2386.174737737738u,0 2386.175737737738u,1.5 2387.1522777777777u,1.5 2387.153277777778u,0 2388.1298178178176u,0 2388.130817817818u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2398.882758258258u,1.5 2398.8837582582582u,0 2400.8378383383383u,0 2400.8388383383385u,1.5 2401.8153783783787u,1.5 2401.816378378379u,0 2402.792918418418u,0 2402.7939184184183u,1.5 2403.7704584584585u,1.5 2403.7714584584587u,0 2405.7255385385383u,0 2405.7265385385385u,1.5 2410.613238738739u,1.5 2410.614238738739u,0 2411.5907787787787u,0 2411.591778778779u,1.5 2412.5683188188186u,1.5 2412.569318818819u,0 2415.500938938939u,0 2415.501938938939u,1.5 2416.478478978979u,1.5 2416.4794789789794u,0 2423.321259259259u,0 2423.322259259259u,1.5 2425.2763393393393u,1.5 2425.2773393393395u,0 2426.2538793793797u,0 2426.25487937938u,1.5 2432.119119619619u,1.5 2432.1201196196193u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2435.05173973974u,0 2435.05273973974u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.9843598598595u,0 2437.9853598598597u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2441.8945200200196u,0 2441.89552002002u,1.5 2442.87206006006u,1.5 2442.87306006006u,0 2446.78222022022u,0 2446.7832202202203u,1.5 2447.75976026026u,1.5 2447.76076026026u,0 2449.7148403403403u,0 2449.7158403403405u,1.5 2451.66992042042u,1.5 2451.6709204204203u,0 2452.6474604604605u,0 2452.6484604604607u,1.5 2454.6025405405403u,1.5 2454.6035405405405u,0 2455.5800805805807u,0 2455.581080580581u,1.5 2459.490240740741u,1.5 2459.491240740741u,0 2462.4228608608605u,0 2462.4238608608607u,1.5 2464.377940940941u,1.5 2464.378940940941u,0 2465.355480980981u,0 2465.3564809809814u,1.5 2466.3330210210206u,1.5 2466.334021021021u,0 2467.310561061061u,0 2467.311561061061u,1.5 2468.288101101101u,1.5 2468.289101101101u,0 2472.198261261261u,0 2472.199261261261u,1.5 2474.1533413413413u,1.5 2474.1543413413415u,0 2476.108421421421u,0 2476.1094214214213u,1.5 2478.0635015015014u,1.5 2478.0645015015016u,0 2482.9512017017014u,0 2482.9522017017016u,1.5 2483.9287417417418u,1.5 2483.929741741742u,0 2484.9062817817817u,0 2484.907281781782u,1.5 2485.8838218218216u,1.5 2485.884821821822u,0 2500.546922422422u,0 2500.5479224224223u,1.5 2505.434622622622u,1.5 2505.4356226226223u,0 2512.277402902903u,0 2512.278402902903u,1.5 2513.2549429429428u,1.5 2513.255942942943u,0 2517.165103103103u,0 2517.166103103103u,1.5 2518.1426431431432u,1.5 2518.1436431431434u,0 2519.120183183183u,0 2519.1211831831833u,1.5 2520.097723223223u,1.5 2520.0987232232233u,0 2522.0528033033033u,0 2522.0538033033035u,1.5 2523.0303433433432u,1.5 2523.0313433433435u,0 2524.985423423423u,0 2524.9864234234233u,1.5 2525.9629634634634u,1.5 2525.9639634634636u,0 2527.9180435435437u,0 2527.919043543544u,1.5 2528.8955835835836u,1.5 2528.896583583584u,0 2529.8731236236235u,0 2529.8741236236237u,1.5 2531.8282037037034u,1.5 2531.8292037037036u,0 2532.8057437437437u,0 2532.806743743744u,1.5 2533.7832837837836u,1.5 2533.784283783784u,0 2534.7608238238236u,0 2534.7618238238238u,1.5 2539.6485240240236u,1.5 2539.649524024024u,0 2540.626064064064u,0 2540.627064064064u,1.5 2544.536224224224u,1.5 2544.5372242242242u,0 2546.4913043043043u,0 2546.4923043043045u,1.5 2547.4688443443442u,1.5 2547.4698443443444u,0 2548.4463843843846u,0 2548.447384384385u,1.5 2549.423924424424u,1.5 2549.4249244244243u,0 2550.4014644644644u,0 2550.4024644644646u,1.5 2552.3565445445447u,1.5 2552.357544544545u,0 2554.3116246246245u,0 2554.3126246246247u,1.5 2556.2667047047044u,1.5 2556.2677047047046u,0 2557.2442447447447u,0 2557.245244744745u,1.5 2562.1319449449447u,1.5 2562.132944944945u,0 2565.064565065065u,0 2565.065565065065u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2567.019645145145u,0 2567.0206451451454u,1.5 2567.997185185185u,1.5 2567.9981851851853u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2577.7725855855856u,1.5 2577.773585585586u,0 2586.5704459459457u,0 2586.571445945946u,1.5 2587.547985985986u,1.5 2587.5489859859863u,0 2588.5255260260255u,0 2588.5265260260257u,1.5 2596.345846346346u,1.5 2596.3468463463464u,0 2597.3233863863866u,0 2597.324386386387u,1.5 2598.300926426426u,1.5 2598.3019264264262u,0 2599.2784664664664u,0 2599.2794664664666u,1.5 2600.2560065065063u,1.5 2600.2570065065065u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2608.0763268268265u,0 2608.0773268268267u,1.5 2611.0089469469467u,1.5 2611.009946946947u,0 2611.986486986987u,0 2611.9874869869873u,1.5 2612.9640270270265u,1.5 2612.9650270270267u,0 2613.941567067067u,0 2613.942567067067u,1.5 2615.896647147147u,1.5 2615.8976471471474u,0 2619.8068073073073u,0 2619.8078073073075u,1.5 2620.784347347347u,1.5 2620.7853473473474u,0 2622.739427427427u,0 2622.740427427427u,1.5 2628.6046676676674u,1.5 2628.6056676676676u,0 2629.5822077077073u,0 2629.5832077077075u,1.5 2630.5597477477477u,1.5 2630.560747747748u,0 2634.469907907908u,0 2634.470907907908u,1.5 2635.4474479479477u,1.5 2635.448447947948u,0 2637.402528028028u,0 2637.403528028028u,1.5 2642.2902282282284u,1.5 2642.2912282282286u,0 2643.267768268268u,0 2643.268768268268u,1.5 2644.2453083083083u,1.5 2644.2463083083085u,0 2651.0880885885886u,0 2651.0890885885888u,1.5 2652.065628628629u,1.5 2652.066628628629u,0 2653.0431686686684u,0 2653.0441686686686u,1.5 2654.9982487487487u,1.5 2654.999248748749u,0 2655.9757887887886u,0 2655.976788788789u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2666.7287292292294u,0 2666.7297292292296u,1.5 2667.706269269269u,1.5 2667.707269269269u,0 2672.5939694694694u,0 2672.5949694694696u,1.5 2673.5715095095093u,1.5 2673.5725095095095u,0 2674.5490495495496u,0 2674.55004954955u,1.5 2679.4367497497497u,1.5 2679.43774974975u,0 2681.39182982983u,0 2681.39282982983u,1.5 2682.3693698698694u,1.5 2682.3703698698696u,0 2684.3244499499497u,0 2684.32544994995u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2689.21215015015u,1.5 2689.2131501501503u,0 2691.1672302302304u,0 2691.1682302302306u,1.5 2693.1223103103102u,1.5 2693.1233103103104u,0 2694.09985035035u,0 2694.1008503503504u,1.5 2695.0773903903905u,1.5 2695.0783903903907u,0 2696.0549304304304u,0 2696.0559304304306u,1.5 2698.0100105105103u,1.5 2698.0110105105105u,0 2698.9875505505506u,0 2698.988550550551u,1.5 2699.9650905905905u,1.5 2699.9660905905907u,0 2701.9201706706704u,0 2701.9211706706706u,1.5 2703.8752507507506u,1.5 2703.876250750751u,0 2706.8078708708704u,0 2706.8088708708706u,1.5 2710.718031031031u,1.5 2710.719031031031u,0 2713.650651151151u,0 2713.6516511511513u,1.5 2714.628191191191u,1.5 2714.6291911911912u,0 2718.538351351351u,0 2718.5393513513513u,1.5 2719.5158913913915u,1.5 2719.5168913913917u,0 2721.4709714714713u,0 2721.4719714714715u,1.5 2722.4485115115112u,1.5 2722.4495115115114u,0 2723.4260515515516u,0 2723.427051551552u,1.5 2725.381131631632u,1.5 2725.382131631632u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2730.268831831832u,0 2730.269831831832u,1.5 2733.2014519519516u,1.5 2733.202451951952u,0 2735.156532032032u,0 2735.157532032032u,1.5 2736.134072072072u,1.5 2736.135072072072u,0 2737.1116121121117u,0 2737.112612112112u,1.5 2738.089152152152u,1.5 2738.0901521521523u,0 2739.066692192192u,0 2739.067692192192u,1.5 2740.0442322322324u,1.5 2740.0452322322326u,0 2741.021772272272u,0 2741.022772272272u,1.5 2745.9094724724723u,1.5 2745.9104724724725u,0 2746.8870125125122u,0 2746.8880125125124u,1.5 2747.8645525525526u,1.5 2747.865552552553u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 2755.6848728728723u,1.5 2755.6858728728726u,0 2756.6624129129127u,0 2756.663412912913u,1.5 2757.6399529529526u,1.5 2757.640952952953u,0 2760.572573073073u,0 2760.573573073073u,1.5 2761.5501131131127u,1.5 2761.551113113113u,0 2762.527653153153u,0 2762.5286531531533u,1.5 2765.460273273273u,1.5 2765.461273273273u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2773.2805935935935u,0 2773.2815935935937u,1.5 2777.1907537537536u,1.5 2777.191753753754u,0 2782.0784539539536u,0 2782.079453953954u,1.5 2786.966154154154u,1.5 2786.9671541541543u,0 2787.943694194194u,0 2787.944694194194u,1.5 2788.9212342342344u,1.5 2788.9222342342346u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2795.764014514514u,1.5 2795.7650145145144u,0 2796.7415545545546u,0 2796.7425545545548u,1.5 2798.696634634635u,1.5 2798.697634634635u,0 2800.6517147147147u,0 2800.652714714715u,1.5 2803.584334834835u,1.5 2803.585334834835u,0 2804.561874874875u,0 2804.562874874875u,1.5 2805.5394149149147u,1.5 2805.540414914915u,0 2806.5169549549546u,0 2806.517954954955u,1.5 2808.472035035035u,1.5 2808.473035035035u,0 2809.449575075075u,0 2809.450575075075u,1.5 2810.4271151151147u,1.5 2810.428115115115u,0 2814.337275275275u,0 2814.338275275275u,1.5 2819.2249754754753u,1.5 2819.2259754754755u,0 2820.202515515515u,0 2820.2035155155154u,1.5 2829.9779159159157u,1.5 2829.978915915916u,0 2831.932995995996u,0 2831.933995995996u,1.5 2833.888076076076u,1.5 2833.889076076076u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2839.753316316316u,1.5 2839.7543163163164u,0 2840.730856356356u,0 2840.7318563563563u,1.5 2844.641016516516u,1.5 2844.6420165165164u,0 2846.5960965965965u,0 2846.5970965965967u,1.5 2847.573636636637u,1.5 2847.574636636637u,0 2848.5511766766763u,0 2848.5521766766765u,1.5 2850.5062567567566u,1.5 2850.5072567567568u,0 2852.461336836837u,0 2852.462336836837u,1.5 2855.3939569569566u,1.5 2855.394956956957u,0 2856.371496996997u,0 2856.372496996997u,1.5 2857.349037037037u,1.5 2857.350037037037u,0 2859.3041171171167u,0 2859.305117117117u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2865.169357357357u,1.5 2865.1703573573573u,0 2866.1468973973974u,0 2866.1478973973976u,1.5 2871.0345975975974u,1.5 2871.0355975975976u,0 2874.9447577577575u,0 2874.9457577577577u,1.5 2876.899837837838u,1.5 2876.900837837838u,0 2877.877377877878u,0 2877.8783778778784u,1.5 2878.8549179179176u,1.5 2878.855917917918u,0 2879.832457957958u,0 2879.833457957958u,1.5 2880.809997997998u,1.5 2880.810997997998u,0 2881.787538038038u,0 2881.788538038038u,1.5 2882.765078078078u,1.5 2882.7660780780784u,0 2883.7426181181177u,0 2883.743618118118u,1.5 2885.697698198198u,1.5 2885.698698198198u,0 2886.6752382382383u,0 2886.6762382382385u,1.5 2887.652778278278u,1.5 2887.6537782782784u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2899.3832587587585u,1.5 2899.3842587587587u,0 2900.360798798799u,0 2900.361798798799u,1.5 2901.338338838839u,1.5 2901.339338838839u,0 2902.315878878879u,0 2902.3168788788794u,1.5 2903.2934189189186u,1.5 2903.294418918919u,0 2909.158659159159u,0 2909.159659159159u,1.5 2910.136199199199u,1.5 2910.137199199199u,0 2912.091279279279u,0 2912.0922792792794u,1.5 2913.068819319319u,1.5 2913.0698193193193u,0 2914.046359359359u,0 2914.0473593593592u,1.5 2921.8666796796797u,1.5 2921.86767967968u,0 2922.8442197197196u,0 2922.84521971972u,1.5 2923.8217597597595u,1.5 2923.8227597597597u,0 2930.66454004004u,0 2930.66554004004u,1.5 2931.64208008008u,1.5 2931.6430800800804u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2938.48486036036u,1.5 2938.48586036036u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 2946.3051806806807u,1.5 2946.306180680681u,0 2947.2827207207206u,0 2947.283720720721u,1.5 2948.2602607607605u,1.5 2948.2612607607607u,0 2949.237800800801u,0 2949.238800800801u,1.5 2950.215340840841u,1.5 2950.216340840841u,0 2955.103041041041u,0 2955.104041041041u,1.5 2956.080581081081u,1.5 2956.0815810810814u,0 2958.035661161161u,0 2958.036661161161u,1.5 2959.013201201201u,1.5 2959.014201201201u,0 2962.923361361361u,0 2962.924361361361u,1.5 2963.9009014014014u,1.5 2963.9019014014016u,0 2965.8559814814816u,0 2965.856981481482u,1.5 2966.833521521521u,1.5 2966.8345215215213u,0 2968.7886016016014u,0 2968.7896016016016u,1.5 2969.7661416416418u,1.5 2969.767141641642u,0 2970.7436816816817u,0 2970.744681681682u,1.5 2971.7212217217216u,1.5 2971.722221721722u,0 2972.6987617617615u,0 2972.6997617617617u,1.5 2973.676301801802u,1.5 2973.677301801802u,0 2974.6538418418418u,0 2974.654841841842u,1.5 2979.541542042042u,1.5 2979.542542042042u,0 2980.519082082082u,0 2980.5200820820824u,1.5 2982.474162162162u,1.5 2982.475162162162u,0 2983.451702202202u,0 2983.452702202202u,1.5 2992.2495625625625u,1.5 2992.2505625625627u,0 2993.2271026026024u,0 2993.2281026026026u,1.5 2999.0923428428428u,1.5 2999.093342842843u,0 3000.069882882883u,0 3000.0708828828833u,1.5 3003.002503003003u,1.5 3003.003503003003u,0 3003.980043043043u,0 3003.9810430430434u,1.5 3006.912663163163u,1.5 3006.913663163163u,0 3009.845283283283u,0 3009.8462832832834u,1.5 3010.822823323323u,1.5 3010.8238233233233u,0 3011.800363363363u,0 3011.801363363363u,1.5 3013.7554434434433u,1.5 3013.7564434434435u,0 3014.7329834834836u,0 3014.733983483484u,1.5 3016.6880635635634u,1.5 3016.6890635635636u,0 3017.6656036036034u,0 3017.6666036036036u,1.5 3018.6431436436437u,1.5 3018.644143643644u,0 3019.6206836836836u,0 3019.621683683684u,1.5 3022.553303803804u,1.5 3022.554303803804u,0 3024.508383883884u,0 3024.5093838838843u,1.5 3025.4859239239236u,1.5 3025.4869239239238u,0 3027.441004004004u,0 3027.442004004004u,1.5 3028.418544044044u,1.5 3028.4195440440444u,0 3029.396084084084u,0 3029.3970840840843u,1.5 3030.373624124124u,1.5 3030.3746241241242u,0 3032.328704204204u,0 3032.329704204204u,1.5 3033.306244244244u,1.5 3033.3072442442444u,0 3034.283784284284u,0 3034.2847842842843u,1.5 3035.261324324324u,1.5 3035.2623243243243u,0 3038.1939444444442u,0 3038.1949444444444u,1.5 3039.1714844844846u,1.5 3039.172484484485u,0 3040.149024524524u,0 3040.1500245245243u,1.5 3041.1265645645644u,1.5 3041.1275645645646u,0 3042.1041046046043u,0 3042.1051046046045u,1.5 3044.0591846846846u,1.5 3044.060184684685u,0 3046.0142647647644u,0 3046.0152647647647u,1.5 3046.991804804805u,1.5 3046.992804804805u,0 3048.946884884885u,0 3048.9478848848853u,1.5 3050.901964964965u,1.5 3050.902964964965u,0 3052.857045045045u,0 3052.8580450450454u,1.5 3054.812125125125u,1.5 3054.813125125125u,0 3055.789665165165u,0 3055.790665165165u,1.5 3062.6324454454452u,1.5 3062.6334454454454u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3066.5426056056053u,0 3066.5436056056055u,1.5 3067.5201456456457u,1.5 3067.521145645646u,0 3073.385385885886u,0 3073.3863858858863u,1.5 3074.3629259259255u,1.5 3074.3639259259257u,0 3077.295546046046u,0 3077.2965460460464u,1.5 3079.250626126126u,1.5 3079.251626126126u,0 3080.228166166166u,0 3080.229166166166u,1.5 3084.138326326326u,1.5 3084.139326326326u,0 3085.115866366366u,0 3085.116866366366u,1.5 3088.0484864864866u,1.5 3088.049486486487u,0 3090.0035665665664u,0 3090.0045665665666u,1.5 3090.9811066066063u,1.5 3090.9821066066065u,0 3092.9361866866866u,0 3092.937186686687u,1.5 3093.9137267267265u,1.5 3093.9147267267267u,0 3094.8912667667664u,0 3094.8922667667666u,1.5 3095.868806806807u,1.5 3095.869806806807u,0 3096.8463468468467u,0 3096.847346846847u,1.5 3097.823886886887u,1.5 3097.8248868868873u,0 3098.8014269269265u,0 3098.8024269269267u,1.5 3102.711587087087u,1.5 3102.7125870870873u,0 3104.666667167167u,0 3104.667667167167u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3112.4869874874876u,0 3112.4879874874878u,1.5 3113.464527527527u,1.5 3113.4655275275272u,0 3114.4420675675674u,0 3114.4430675675676u,1.5 3115.4196076076073u,1.5 3115.4206076076075u,0 3116.3971476476477u,0 3116.398147647648u,1.5 3118.3522277277275u,1.5 3118.3532277277277u,0 3120.307307807808u,0 3120.308307807808u,1.5 3122.262387887888u,1.5 3122.2633878878883u,0 3125.195008008008u,0 3125.196008008008u,1.5 3126.172548048048u,1.5 3126.1735480480484u,0 3127.150088088088u,0 3127.1510880880883u,1.5 3128.127628128128u,1.5 3128.128628128128u,0 3131.060248248248u,0 3131.0612482482484u,1.5 3135.947948448448u,1.5 3135.9489484484484u,0 3139.8581086086083u,0 3139.8591086086085u,1.5 3140.8356486486487u,1.5 3140.836648648649u,0 3143.7682687687684u,0 3143.7692687687686u,1.5 3147.678428928929u,1.5 3147.679428928929u,0 3148.655968968969u,0 3148.656968968969u,1.5 3151.588589089089u,1.5 3151.5895890890893u,0 3153.543669169169u,0 3153.544669169169u,1.5 3154.5212092092092u,1.5 3154.5222092092094u,0 3155.498749249249u,0 3155.4997492492494u,1.5 3156.476289289289u,1.5 3156.4772892892893u,0 3157.4538293293294u,0 3157.4548293293296u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3168.2067697697694u,0 3168.2077697697696u,1.5 3169.1843098098097u,1.5 3169.18530980981u,0 3170.1618498498497u,0 3170.16284984985u,1.5 3175.04955005005u,1.5 3175.0505500500503u,0 3177.0046301301304u,0 3177.0056301301306u,1.5 3178.9597102102102u,1.5 3178.9607102102104u,0 3179.93725025025u,0 3179.9382502502503u,1.5 3180.91479029029u,1.5 3180.9157902902903u,0 3182.86987037037u,0 3182.87087037037u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3190.6901906906905u,0 3190.6911906906907u,1.5 3191.667730730731u,1.5 3191.668730730731u,0 3192.6452707707704u,0 3192.6462707707706u,1.5 3196.555430930931u,1.5 3196.556430930931u,0 3197.532970970971u,0 3197.533970970971u,1.5 3198.5105110110107u,1.5 3198.511511011011u,0 3202.420671171171u,0 3202.421671171171u,1.5 3203.398211211211u,1.5 3203.3992112112114u,0 3204.375751251251u,0 3204.3767512512513u,1.5 3207.308371371371u,1.5 3207.309371371371u,0 3213.1736116116112u,0 3213.1746116116115u,1.5 3215.1286916916915u,1.5 3215.1296916916917u,0 3217.0837717717714u,0 3217.0847717717716u,1.5 3218.0613118118117u,1.5 3218.062311811812u,0 3219.0388518518516u,0 3219.039851851852u,1.5 3220.016391891892u,1.5 3220.017391891892u,0 3223.926552052052u,0 3223.9275520520523u,1.5 3224.904092092092u,1.5 3224.905092092092u,0 3225.8816321321324u,0 3225.8826321321326u,1.5 3227.836712212212u,1.5 3227.8377122122124u,0 3228.814252252252u,0 3228.8152522522523u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3232.724412412412u,0 3232.7254124124124u,1.5 3234.6794924924925u,1.5 3234.6804924924927u,0 3236.6345725725723u,0 3236.6355725725725u,1.5 3237.6121126126122u,1.5 3237.6131126126124u,0 3238.5896526526526u,0 3238.590652652653u,1.5 3239.5671926926925u,1.5 3239.5681926926927u,0 3240.544732732733u,0 3240.545732732733u,1.5 3242.4998128128127u,1.5 3242.500812812813u,0 3244.454892892893u,0 3244.455892892893u,1.5 3245.432432932933u,1.5 3245.433432932933u,0 3246.409972972973u,0 3246.410972972973u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3255.2078333333334u,0 3255.2088333333336u,1.5 3259.1179934934935u,1.5 3259.1189934934937u,0 3260.0955335335334u,0 3260.0965335335336u,1.5 3262.050613613613u,1.5 3262.0516136136134u,0 3263.0281536536536u,0 3263.029153653654u,1.5 3264.0056936936935u,1.5 3264.0066936936937u,0 3264.983233733734u,0 3264.984233733734u,1.5 3265.9607737737733u,1.5 3265.9617737737735u,0 3267.9158538538536u,0 3267.916853853854u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3274.7586341341344u,1.5 3274.7596341341346u,0 3277.691254254254u,0 3277.6922542542543u,1.5 3278.6687942942945u,1.5 3278.6697942942947u,0 3279.6463343343344u,0 3279.6473343343346u,1.5 3280.6238743743743u,1.5 3280.6248743743745u,0 3281.601414414414u,0 3281.6024144144144u,1.5 3283.5564944944945u,1.5 3283.5574944944947u,0 3285.5115745745743u,0 3285.5125745745745u,1.5 3286.489114614614u,1.5 3286.4901146146144u,0 3287.4666546546546u,0 3287.467654654655u,1.5 3289.421734734735u,1.5 3289.422734734735u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3294.309434934935u,1.5 3294.310434934935u,0 3297.242055055055u,0 3297.2430550550553u,1.5 3298.219595095095u,1.5 3298.220595095095u,0 3299.1971351351353u,0 3299.1981351351355u,1.5 3302.129755255255u,1.5 3302.1307552552553u,0 3303.1072952952954u,0 3303.1082952952956u,1.5 3304.0848353353354u,1.5 3304.0858353353356u,0 3307.9949954954955u,0 3307.9959954954957u,1.5 3308.9725355355354u,1.5 3308.9735355355356u,0 3310.927615615615u,0 3310.9286156156154u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3320.7030160160157u,0 3320.704016016016u,1.5 3325.590716216216u,1.5 3325.5917162162164u,0 3330.478416416416u,0 3330.4794164164164u,1.5 3331.455956456456u,1.5 3331.4569564564563u,0 3332.4334964964964u,0 3332.4344964964966u,1.5 3334.3885765765763u,1.5 3334.3895765765765u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3345.1415170170167u,0 3345.142517017017u,1.5 3347.096597097097u,1.5 3347.097597097097u,0 3348.0741371371373u,0 3348.0751371371375u,1.5 3349.0516771771768u,1.5 3349.052677177177u,0 3350.029217217217u,0 3350.0302172172173u,1.5 3351.006757257257u,1.5 3351.0077572572573u,0 3351.9842972972974u,0 3351.9852972972976u,1.5 3352.9618373373373u,1.5 3352.9628373373375u,0 3353.9393773773772u,0 3353.9403773773774u,1.5 3355.894457457457u,1.5 3355.8954574574573u,0 3357.8495375375373u,0 3357.8505375375375u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3365.6698578578576u,0 3365.6708578578578u,1.5 3366.647397897898u,1.5 3366.648397897898u,0 3369.5800180180177u,0 3369.581018018018u,1.5 3370.557558058058u,1.5 3370.558558058058u,0 3371.535098098098u,0 3371.536098098098u,1.5 3378.3778783783787u,1.5 3378.378878378379u,0 3382.2880385385383u,0 3382.2890385385385u,1.5 3384.243118618618u,1.5 3384.2441186186184u,0 3385.2206586586585u,0 3385.2216586586587u,1.5 3386.1981986986984u,1.5 3386.1991986986986u,0 3387.175738738739u,0 3387.176738738739u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3390.1083588588585u,0 3390.1093588588587u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.996059059059u,0 3394.997059059059u,1.5 3396.9511391391393u,1.5 3396.9521391391395u,0 3401.8388393393393u,0 3401.8398393393395u,1.5 3402.8163793793797u,1.5 3402.81737937938u,0 3404.7714594594595u,0 3404.7724594594597u,1.5 3409.6591596596595u,1.5 3409.6601596596597u,0 3410.6366996996994u,0 3410.6376996996996u,1.5 3413.5693198198196u,1.5 3413.57031981982u,0 3414.5468598598595u,0 3414.5478598598597u,1.5 3419.43456006006u,1.5 3419.43556006006u,0 3420.4121001001u,0 3420.4131001001u,1.5 3421.3896401401403u,1.5 3421.3906401401405u,0 3422.36718018018u,0 3422.3681801801804u,1.5 3423.34472022022u,1.5 3423.3457202202203u,0 3424.32226026026u,0 3424.32326026026u,1.5 3426.2773403403403u,1.5 3426.2783403403405u,0 3427.2548803803807u,0 3427.255880380381u,1.5 3430.1875005005004u,1.5 3430.1885005005006u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3434.0976606606605u,1.5 3434.0986606606607u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3436.052740740741u,1.5 3436.053740740741u,0 3450.7158413413413u,0 3450.7168413413415u,1.5 3451.6933813813816u,1.5 3451.694381381382u,0 3452.670921421421u,0 3452.6719214214213u,1.5 3454.6260015015014u,1.5 3454.6270015015016u,0 3457.558621621621u,0 3457.5596216216213u,1.5 3458.5361616616615u,1.5 3458.5371616616617u,0 3459.5137017017014u,0 3459.5147017017016u,1.5 3463.4238618618615u,1.5 3463.4248618618617u,0 3464.401401901902u,0 3464.402401901902u,1.5 3466.356481981982u,1.5 3466.3574819819823u,0 3468.311562062062u,0 3468.312562062062u,1.5 3469.289102102102u,1.5 3469.290102102102u,0 3471.244182182182u,0 3471.2451821821824u,1.5 3472.221722222222u,1.5 3472.2227222222223u,0 3475.1543423423423u,0 3475.1553423423425u,1.5 3476.1318823823826u,1.5 3476.132882382383u,0 3478.0869624624625u,0 3478.0879624624627u,1.5 3480.0420425425427u,1.5 3480.043042542543u,0 3484.9297427427427u,0 3484.930742742743u,1.5 3485.9072827827827u,1.5 3485.908282782783u,0 3486.8848228228226u,0 3486.885822822823u,1.5 3489.8174429429428u,1.5 3489.818442942943u,0 3494.7051431431432u,0 3494.7061431431434u,1.5 3495.682683183183u,1.5 3495.6836831831833u,0 3496.660223223223u,0 3496.6612232232233u,1.5 3498.6153033033033u,1.5 3498.6163033033035u,0 3500.5703833833836u,0 3500.571383383384u,1.5 3501.547923423423u,1.5 3501.5489234234233u,0 3511.3233238238236u,0 3511.3243238238238u,1.5 3512.3008638638635u,1.5 3512.3018638638637u,0 3513.278403903904u,0 3513.279403903904u,1.5 3515.233483983984u,1.5 3515.2344839839843u,0 3521.098724224224u,0 3521.0997242242242u,1.5 3522.076264264264u,1.5 3522.077264264264u,0 3524.0313443443442u,0 3524.0323443443444u,1.5 3525.986424424424u,1.5 3525.9874244244243u,0 3527.9415045045043u,0 3527.9425045045045u,1.5 3528.9190445445447u,1.5 3528.920044544545u,0 3529.8965845845846u,0 3529.897584584585u,1.5 3530.8741246246245u,1.5 3530.8751246246247u,0 3532.8292047047044u,0 3532.8302047047046u,1.5 3538.6944449449447u,1.5 3538.695444944945u,0 3539.671984984985u,0 3539.6729849849853u,1.5 3544.559685185185u,1.5 3544.5606851851853u,0 3545.537225225225u,0 3545.5382252252252u,1.5 3549.4473853853856u,1.5 3549.448385385386u,0 3551.4024654654654u,0 3551.4034654654656u,1.5 3552.3800055055053u,1.5 3552.3810055055055u,0 3553.3575455455457u,0 3553.358545545546u,1.5 3554.3350855855856u,1.5 3554.336085585586u,0 3556.2901656656654u,0 3556.2911656656656u,1.5 3557.2677057057053u,1.5 3557.2687057057055u,0 3562.155405905906u,0 3562.156405905906u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.020646146146u,1.5 3568.0216461461464u,0 3569.975726226226u,0 3569.976726226226u,1.5 3571.9308063063063u,1.5 3571.9318063063065u,0 3572.908346346346u,0 3572.9093463463464u,1.5 3574.863426426426u,1.5 3574.8644264264262u,0 3576.8185065065063u,0 3576.8195065065065u,1.5 3579.7511266266265u,1.5 3579.7521266266267u,0 3586.593906906907u,0 3586.594906906907u,1.5 3587.5714469469467u,1.5 3587.572446946947u,0 3588.548986986987u,0 3588.5499869869873u,1.5 3591.481607107107u,1.5 3591.482607107107u,0 3592.459147147147u,0 3592.4601471471474u,1.5 3593.436687187187u,1.5 3593.4376871871873u,0 3594.414227227227u,0 3594.415227227227u,1.5 3595.391767267267u,1.5 3595.392767267267u,0 3596.3693073073073u,0 3596.3703073073075u,1.5 3597.346847347347u,1.5 3597.3478473473474u,0 3598.3243873873876u,0 3598.3253873873878u,1.5 3599.301927427427u,1.5 3599.302927427427u,0 3602.2345475475477u,0 3602.235547547548u,1.5 3605.1671676676674u,1.5 3605.1681676676676u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3607.1222477477477u,1.5 3607.123247747748u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3612.987487987988u,1.5 3612.9884879879883u,0 3613.9650280280275u,0 3613.9660280280277u,1.5 3614.942568068068u,1.5 3614.943568068068u,0 3621.785348348348u,0 3621.7863483483484u,1.5 3623.740428428428u,1.5 3623.741428428428u,0 3624.7179684684684u,0 3624.7189684684686u,1.5 3629.6056686686684u,1.5 3629.6066686686686u,0 3635.4709089089088u,0 3635.471908908909u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3637.425988988989u,0 3637.4269889889893u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3640.358609109109u,1.5 3640.359609109109u,0 3641.336149149149u,0 3641.3371491491494u,1.5 3644.268769269269u,1.5 3644.269769269269u,0 3645.2463093093093u,0 3645.2473093093095u,1.5 3647.2013893893895u,1.5 3647.2023893893897u,0 3651.1115495495496u,0 3651.11254954955u,1.5 3653.06662962963u,1.5 3653.06762962963u,0 3654.0441696696694u,0 3654.0451696696696u,1.5 3655.0217097097097u,1.5 3655.02270970971u,0 3656.9767897897896u,0 3656.9777897897898u,1.5 3657.95432982983u,1.5 3657.95532982983u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3669.6848103103102u,1.5 3669.6858103103104u,0 3673.5949704704703u,0 3673.5959704704705u,1.5 3674.5725105105103u,1.5 3674.5735105105105u,0 3675.5500505505506u,0 3675.551050550551u,1.5 3678.4826706706704u,1.5 3678.4836706706706u,0 3679.4602107107107u,0 3679.461210710711u,1.5 3680.4377507507506u,1.5 3680.438750750751u,0 3681.4152907907906u,0 3681.4162907907908u,1.5 3682.392830830831u,1.5 3682.393830830831u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3689.2356111111108u,0 3689.236611111111u,1.5 3690.213151151151u,1.5 3690.2141511511513u,0 3691.190691191191u,0 3691.1916911911912u,1.5 3693.145771271271u,1.5 3693.146771271271u,0 3697.0559314314314u,0 3697.0569314314316u,1.5 3699.9885515515516u,1.5 3699.989551551552u,0 3700.9660915915915u,0 3700.9670915915917u,1.5 3702.9211716716713u,1.5 3702.9221716716715u,0 3706.831331831832u,0 3706.832331831832u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3711.719032032032u,1.5 3711.720032032032u,0 3715.629192192192u,0 3715.630192192192u,1.5 3716.6067322322324u,1.5 3716.6077322322326u,0 3717.584272272272u,0 3717.585272272272u,1.5 3719.539352352352u,1.5 3719.5403523523523u,0 3722.4719724724723u,0 3722.4729724724725u,1.5 3723.4495125125122u,1.5 3723.4505125125124u,0 3724.4270525525526u,0 3724.428052552553u,1.5 3725.4045925925925u,1.5 3725.4055925925927u,0 3730.292292792793u,0 3730.293292792793u,1.5 3732.2473728728723u,1.5 3732.2483728728726u,0 3734.2024529529526u,0 3734.203452952953u,1.5 3735.179992992993u,1.5 3735.180992992993u,0 3736.157533033033u,0 3736.158533033033u,1.5 3737.135073073073u,1.5 3737.136073073073u,0 3739.090153153153u,0 3739.0911531531533u,1.5 3740.067693193193u,1.5 3740.068693193193u,0 3741.0452332332334u,0 3741.0462332332336u,1.5 3744.9553933933935u,1.5 3744.9563933933937u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3753.7532537537536u,0 3753.754253753754u,1.5 3754.730793793794u,1.5 3754.731793793794u,0 3755.708333833834u,0 3755.709333833834u,1.5 3756.685873873874u,1.5 3756.686873873874u,0 3757.6634139139137u,0 3757.664413913914u,1.5 3758.6409539539536u,1.5 3758.641953953954u,0 3759.618493993994u,0 3759.619493993994u,1.5 3760.596034034034u,1.5 3760.597034034034u,0 3761.573574074074u,0 3761.574574074074u,1.5 3764.506194194194u,1.5 3764.507194194194u,0 3772.326514514514u,0 3772.3275145145144u,1.5 3774.2815945945945u,1.5 3774.2825945945947u,0 3775.259134634635u,0 3775.260134634635u,1.5 3776.2366746746743u,1.5 3776.2376746746745u,0 3778.1917547547546u,0 3778.192754754755u,1.5 3779.169294794795u,1.5 3779.170294794795u,0 3780.146834834835u,0 3780.147834834835u,1.5 3781.124374874875u,1.5 3781.125374874875u,0 3783.0794549549546u,0 3783.080454954955u,1.5 3786.012075075075u,1.5 3786.013075075075u,0 3787.967155155155u,0 3787.9681551551553u,1.5 3788.944695195195u,1.5 3788.945695195195u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3793.8323953953955u,1.5 3793.8333953953957u,0 3794.8099354354354u,0 3794.8109354354356u,1.5 3798.7200955955955u,1.5 3798.7210955955957u,0 3802.6302557557556u,0 3802.631255755756u,1.5 3803.607795795796u,1.5 3803.608795795796u,0 3804.585335835836u,0 3804.586335835836u,1.5 3806.5404159159157u,1.5 3806.541415915916u,0 3808.495495995996u,0 3808.496495995996u,1.5 3809.473036036036u,1.5 3809.474036036036u,0 3812.405656156156u,0 3812.4066561561563u,1.5 3813.383196196196u,1.5 3813.384196196196u,0 3814.3607362362363u,0 3814.3617362362365u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3821.203516516516u,0 3821.2045165165164u,1.5 3822.1810565565565u,1.5 3822.1820565565567u,0 3825.1136766766763u,0 3825.1146766766765u,1.5 3826.0912167167166u,1.5 3826.092216716717u,0 3828.046296796797u,0 3828.047296796797u,1.5 3831.9564569569566u,1.5 3831.957456956957u,0 3832.933996996997u,0 3832.934996996997u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3836.844157157157u,1.5 3836.8451571571572u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 3844.6644774774772u,1.5 3844.6654774774775u,0 3847.5970975975974u,0 3847.5980975975976u,1.5 3848.574637637638u,1.5 3848.575637637638u,0 3850.5297177177176u,0 3850.530717717718u,1.5 3851.5072577577575u,1.5 3851.5082577577577u,0 3852.484797797798u,0 3852.485797797798u,1.5 3855.4174179179176u,1.5 3855.418417917918u,0 3856.394957957958u,0 3856.395957957958u,1.5 3859.3275780780777u,1.5 3859.328578078078u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3870.080518518518u,1.5 3870.0815185185184u,0 3873.013138638639u,0 3873.014138638639u,1.5 3873.9906786786783u,1.5 3873.9916786786785u,0 3876.923298798799u,0 3876.924298798799u,1.5 3877.900838838839u,1.5 3877.901838838839u,0 3879.8559189189186u,0 3879.856918918919u,1.5 3888.653779279279u,1.5 3888.6547792792794u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3895.4965595595595u,0 3895.4975595595597u,1.5 3902.33933983984u,1.5 3902.34033983984u,0 3903.31687987988u,0 3903.3178798798804u,1.5 3904.2944199199196u,1.5 3904.29541991992u,0 3913.09228028028u,0 3913.0932802802804u,1.5 3914.06982032032u,1.5 3914.0708203203203u,0 3915.0473603603605u,0 3915.0483603603607u,1.5 3917.00244044044u,1.5 3917.00344044044u,0 3917.9799804804807u,0 3917.980980480481u,1.5 3919.935060560561u,1.5 3919.936060560561u,0 3920.9126006006004u,0 3920.9136006006006u,1.5 3923.8452207207206u,1.5 3923.846220720721u,0 3925.800300800801u,0 3925.801300800801u,1.5 3926.7778408408403u,1.5 3926.7788408408405u,0 3928.7329209209206u,0 3928.733920920921u,1.5 3929.710460960961u,1.5 3929.711460960961u,0 3933.6206211211206u,0 3933.621621121121u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3938.508321321321u,1.5 3938.5093213213213u,0 3939.4858613613615u,0 3939.4868613613617u,1.5 3940.4634014014014u,1.5 3940.4644014014016u,0 3941.440941441441u,0 3941.441941441441u,1.5 3943.396021521521u,1.5 3943.3970215215213u,0 3944.373561561562u,0 3944.374561561562u,1.5 3947.3061816816817u,1.5 3947.307181681682u,0 3948.2837217217216u,0 3948.284721721722u,1.5 3949.261261761762u,1.5 3949.262261761762u,0 3950.238801801802u,0 3950.239801801802u,1.5 3952.193881881882u,1.5 3952.1948818818823u,0 3953.1714219219216u,0 3953.172421921922u,1.5 3954.1489619619624u,1.5 3954.1499619619626u,0 3956.104042042042u,0 3956.105042042042u,1.5 3957.081582082082u,1.5 3957.0825820820824u,0 3960.014202202202u,0 3960.015202202202u,1.5 3961.969282282282u,1.5 3961.9702822822824u,0 3962.946822322322u,0 3962.9478223223223u,1.5 3963.9243623623624u,1.5 3963.9253623623626u,0 3965.879442442442u,0 3965.880442442442u,1.5 3966.8569824824826u,1.5 3966.857982482483u,0 3967.834522522522u,0 3967.8355225225223u,1.5 3969.7896026026024u,1.5 3969.7906026026026u,0 3972.7222227227226u,0 3972.7232227227228u,1.5 3973.699762762763u,1.5 3973.700762762763u,0 3974.677302802803u,0 3974.678302802803u,1.5 3975.6548428428423u,1.5 3975.6558428428425u,0 3977.6099229229226u,0 3977.610922922923u,1.5 3980.5425430430428u,1.5 3980.543543043043u,0 3981.520083083083u,0 3981.5210830830833u,1.5 3982.4976231231226u,1.5 3982.498623123123u,0 3983.4751631631634u,0 3983.4761631631636u,1.5 3989.3404034034033u,1.5 3989.3414034034035u,0 3991.2954834834836u,0 3991.296483483484u,1.5 3998.138263763764u,1.5 3998.139263763764u,0 3999.115803803804u,0 3999.116803803804u,1.5 4000.0933438438433u,1.5 4000.0943438438435u,0 4001.070883883884u,0 4001.0718838838843u,1.5 4013.7789044044043u,1.5 4013.7799044044045u,0 4014.756444444444u,0 4014.757444444444u,1.5 4016.711524524524u,1.5 4016.7125245245243u,0 4018.6666046046043u,0 4018.6676046046045u,1.5 4020.6216846846846u,1.5 4020.622684684685u,0 4021.5992247247245u,0 4021.6002247247247u,1.5 4024.5318448448443u,1.5 4024.5328448448445u,0 4026.4869249249246u,0 4026.4879249249248u,1.5 4027.4644649649654u,1.5 4027.4654649649656u,0 4028.442005005005u,0 4028.443005005005u,1.5 4029.4195450450447u,1.5 4029.420545045045u,0 4030.397085085085u,0 4030.3980850850853u,1.5 4031.374625125125u,1.5 4031.375625125125u,0 4033.329705205205u,0 4033.330705205205u,1.5 4035.284785285285u,1.5 4035.2857852852853u,0 4037.2398653653654u,0 4037.2408653653656u,1.5 4038.2174054054053u,1.5 4038.2184054054055u,0 4039.194945445445u,0 4039.195945445445u,1.5 4040.1724854854856u,1.5 4040.173485485486u,0 4043.1051056056053u,0 4043.1061056056055u,1.5 4045.0601856856856u,1.5 4045.061185685686u,0 4047.015265765766u,0 4047.016265765766u,1.5 4048.9703458458453u,1.5 4048.9713458458455u,0 4049.947885885886u,0 4049.9488858858863u,1.5 4051.9029659659664u,1.5 4051.9039659659666u,0 4052.880506006006u,0 4052.881506006006u,1.5 4057.768206206206u,1.5 4057.769206206206u,0 4058.7457462462457u,0 4058.746746246246u,1.5 4061.6783663663664u,1.5 4061.6793663663666u,0 4062.6559064064063u,0 4062.6569064064065u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4065.588526526526u,0 4065.5895265265262u,1.5 4066.566066566567u,1.5 4066.567066566567u,0 4067.5436066066063u,0 4067.5446066066065u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4073.4088468468462u,0 4073.4098468468464u,1.5 4074.386386886887u,1.5 4074.3873868868873u,0 4075.3639269269265u,0 4075.3649269269267u,1.5 4076.3414669669673u,1.5 4076.3424669669675u,0 4077.319007007007u,0 4077.320007007007u,1.5 4078.2965470470467u,1.5 4078.297547047047u,0 4079.274087087087u,0 4079.2750870870873u,1.5 4080.251627127127u,1.5 4080.252627127127u,0 4081.2291671671674u,0 4081.2301671671676u,1.5 4084.161787287287u,1.5 4084.1627872872873u,0 4085.139327327327u,0 4085.140327327327u,1.5 4086.1168673673674u,1.5 4086.1178673673676u,0 4087.0944074074073u,0 4087.0954074074075u,1.5 4089.0494874874876u,1.5 4089.0504874874878u,0 4092.959647647647u,0 4092.9606476476474u,1.5 4095.892267767768u,1.5 4095.893267767768u,0 4096.869807807808u,0 4096.870807807808u,1.5 4097.847347847847u,1.5 4097.848347847847u,0 4098.824887887888u,0 4098.825887887888u,1.5 4101.757508008008u,1.5 4101.758508008008u,0 4102.735048048047u,0 4102.736048048047u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4105.667668168168u,0 4105.668668168169u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4112.510448448448u,0 4112.511448448448u,1.5 4113.487988488489u,1.5 4113.488988488489u,0 4114.465528528528u,0 4114.466528528528u,1.5 4115.443068568568u,1.5 4115.444068568569u,0 4116.420608608609u,0 4116.421608608609u,1.5 4119.353228728728u,1.5 4119.354228728728u,0 4120.330768768769u,0 4120.3317687687695u,1.5 4122.285848848848u,1.5 4122.286848848848u,0 4124.240928928929u,0 4124.241928928929u,1.5 4125.218468968969u,1.5 4125.2194689689695u,0 4127.173549049048u,0 4127.174549049048u,1.5 4128.1510890890895u,1.5 4128.15208908909u,0 4130.106169169169u,0 4130.1071691691695u,1.5 4131.083709209209u,1.5 4131.084709209209u,0 4132.061249249249u,0 4132.062249249249u,1.5 4134.993869369369u,1.5 4134.99486936937u,0 4137.9264894894895u,0 4137.92748948949u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4140.85910960961u,0 4140.86010960961u,1.5 4141.836649649649u,1.5 4141.837649649649u,0 4142.81418968969u,0 4142.81518968969u,1.5 4144.76926976977u,1.5 4144.7702697697705u,0 4145.74680980981u,0 4145.74780980981u,1.5 4146.724349849849u,1.5 4146.725349849849u,0 4149.65696996997u,0 4149.6579699699705u,1.5 4150.63451001001u,1.5 4150.63551001001u,0 4154.54467017017u,0 4154.5456701701705u,1.5 4155.52221021021u,1.5 4155.52321021021u,0 4156.49975025025u,0 4156.50075025025u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4166.27515065065u,0 4166.27615065065u,1.5 4167.2526906906905u,1.5 4167.253690690691u,0 4168.23023073073u,0 4168.23123073073u,1.5 4170.185310810811u,1.5 4170.186310810811u,0 4171.16285085085u,0 4171.16385085085u,1.5 4172.140390890891u,1.5 4172.141390890891u,0 4173.117930930931u,0 4173.118930930931u,1.5 4174.095470970971u,1.5 4174.0964709709715u,0 4178.005631131131u,0 4178.006631131131u,1.5 4178.983171171171u,1.5 4178.9841711711715u,0 4179.960711211211u,0 4179.961711211211u,1.5 4182.893331331331u,1.5 4182.894331331331u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4190.713651651651u,0 4190.714651651651u,1.5 4192.668731731731u,1.5 4192.669731731731u,0 4194.623811811812u,0 4194.624811811812u,1.5 4197.556431931932u,1.5 4197.557431931932u,0 4198.533971971972u,0 4198.5349719719725u,1.5 4199.511512012012u,1.5 4199.512512012012u,0 4201.4665920920925u,0 4201.467592092093u,1.5 4202.444132132132u,1.5 4202.445132132132u,0 4203.421672172172u,0 4203.4226721721725u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4210.264452452452u,1.5 4210.265452452452u,0 4213.197072572572u,0 4213.1980725725725u,1.5 4216.1296926926925u,1.5 4216.130692692693u,0 4217.107232732732u,0 4217.108232732732u,1.5 4219.062312812813u,1.5 4219.063312812813u,0 4222.972472972973u,0 4222.9734729729735u,1.5 4223.950013013013u,1.5 4223.951013013013u,0 4226.882633133133u,0 4226.883633133133u,1.5 4229.815253253253u,1.5 4229.816253253253u,0 4234.702953453453u,0 4234.703953453453u,1.5 4236.658033533533u,1.5 4236.659033533533u,0 4239.590653653653u,0 4239.591653653653u,1.5 4240.5681936936935u,1.5 4240.569193693694u,0 4244.478353853853u,0 4244.479353853853u,1.5 4245.4558938938935u,1.5 4245.456893893894u,0 4246.433433933934u,0 4246.434433933934u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4254.253754254254u,0 4254.254754254254u,1.5 4255.2312942942945u,1.5 4255.232294294295u,0 4256.208834334334u,0 4256.209834334334u,1.5 4260.1189944944945u,1.5 4260.119994494495u,0 4261.096534534534u,0 4261.097534534534u,1.5 4262.074074574574u,1.5 4262.0750745745745u,0 4265.0066946946945u,0 4265.007694694695u,1.5 4266.961774774775u,1.5 4266.962774774775u,0 4267.939314814815u,0 4267.940314814815u,1.5 4268.916854854855u,1.5 4268.917854854855u,0 4270.871934934935u,0 4270.872934934935u,1.5 4272.827015015015u,1.5 4272.828015015015u,0 4274.782095095095u,0 4274.783095095096u,1.5 4275.759635135135u,1.5 4275.760635135135u,0 4276.737175175175u,0 4276.7381751751755u,1.5 4277.714715215215u,1.5 4277.715715215215u,0 4278.692255255256u,0 4278.693255255256u,1.5 4282.602415415415u,1.5 4282.603415415415u,0 4285.535035535535u,0 4285.536035535535u,1.5 4286.512575575575u,1.5 4286.5135755755755u,0 4288.467655655656u,0 4288.468655655656u,1.5 4289.4451956956955u,1.5 4289.446195695696u,0 4290.422735735735u,0 4290.423735735735u,1.5 4292.377815815816u,1.5 4292.378815815816u,0 4293.355355855856u,0 4293.356355855856u,1.5 4294.3328958958955u,1.5 4294.333895895896u,0 4298.243056056056u,0 4298.244056056056u,1.5 4299.220596096096u,1.5 4299.221596096097u,0 4300.198136136136u,0 4300.199136136136u,1.5 4303.130756256257u,1.5 4303.131756256257u,0 4307.040916416417u,0 4307.041916416417u,1.5 4308.018456456457u,1.5 4308.019456456457u,0 4308.995996496496u,0 4308.996996496497u,1.5 4309.973536536536u,1.5 4309.974536536536u,0 4310.951076576576u,0 4310.9520765765765u,1.5 4313.8836966966965u,1.5 4313.884696696697u,0 4317.793856856857u,0 4317.794856856857u,1.5 4318.7713968968965u,1.5 4318.772396896897u,0 4320.726476976977u,0 4320.727476976977u,1.5 4321.704017017017u,1.5 4321.705017017017u,0 4323.659097097097u,0 4323.660097097098u,1.5 4326.591717217217u,1.5 4326.592717217217u,0 4327.569257257258u,0 4327.570257257258u,1.5 4328.546797297297u,1.5 4328.547797297298u,0 4332.456957457458u,0 4332.457957457458u,1.5 4336.367117617618u,1.5 4336.368117617618u,0 4337.344657657658u,0 4337.345657657658u,1.5 4343.2098978978975u,1.5 4343.210897897898u,0 4344.187437937938u,0 4344.188437937938u,1.5 4345.164977977978u,1.5 4345.165977977978u,0 4346.142518018018u,0 4346.143518018018u,1.5 4347.120058058058u,1.5 4347.121058058058u,0 4348.097598098098u,0 4348.098598098099u,1.5 4351.030218218218u,1.5 4351.031218218218u,0 4354.940378378378u,0 4354.941378378378u,1.5 4355.917918418419u,1.5 4355.918918418419u,0 4357.872998498498u,0 4357.873998498499u,1.5 4358.850538538538u,1.5 4358.851538538538u,0 4359.828078578578u,0 4359.829078578578u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4362.760698698698u,0 4362.761698698699u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4368.625938938939u,0 4368.626938938939u,1.5 4370.581019019019u,1.5 4370.582019019019u,0 4371.558559059059u,0 4371.559559059059u,1.5 4372.536099099099u,1.5 4372.5370990991u,0 4374.491179179179u,0 4374.492179179179u,1.5 4375.468719219219u,1.5 4375.469719219219u,0 4377.423799299299u,0 4377.4247992993u,1.5 4379.378879379379u,1.5 4379.379879379379u,0 4382.311499499499u,0 4382.3124994995u,1.5 4383.289039539539u,1.5 4383.290039539539u,0 4385.24411961962u,0 4385.24511961962u,1.5 4386.22165965966u,1.5 4386.22265965966u,0 4387.199199699699u,0 4387.2001996997u,1.5 4390.13181981982u,1.5 4390.13281981982u,0 4391.10935985986u,0 4391.11035985986u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.99706006006u,1.5 4395.99806006006u,0 4402.83984034034u,0 4402.84084034034u,1.5 4403.81738038038u,1.5 4403.81838038038u,0 4404.794920420421u,0 4404.795920420421u,1.5 4405.772460460461u,1.5 4405.773460460461u,0 4406.7500005005u,0 4406.751000500501u,1.5 4411.6377007007u,1.5 4411.638700700701u,0 4412.61524074074u,0 4412.61624074074u,1.5 4414.570320820821u,1.5 4414.571320820821u,0 4416.5254009009u,0 4416.526400900901u,1.5 4417.502940940941u,1.5 4417.503940940941u,0 4418.480480980981u,0 4418.481480980981u,1.5 4419.458021021021u,1.5 4419.459021021021u,0 4420.435561061061u,0 4420.436561061061u,1.5 4421.413101101101u,1.5 4421.414101101102u,0 4423.368181181181u,0 4423.369181181181u,1.5 4424.345721221221u,1.5 4424.346721221221u,0 4425.323261261262u,0 4425.324261261262u,1.5 4426.300801301301u,1.5 4426.301801301302u,0 4427.278341341341u,0 4427.279341341341u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4438.031281781782u,1.5 4438.032281781782u,0 4440.963901901901u,0 4440.964901901902u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4442.918981981982u,0 4442.919981981982u,1.5 4443.896522022022u,1.5 4443.897522022022u,0 4448.784222222222u,0 4448.785222222222u,1.5 4450.739302302302u,1.5 4450.740302302303u,0 4451.716842342342u,0 4451.717842342342u,1.5 4452.694382382382u,1.5 4452.695382382382u,0 4453.6719224224225u,0 4453.672922422423u,1.5 4456.604542542542u,1.5 4456.605542542542u,0 4457.582082582582u,0 4457.583082582582u,1.5 4459.537162662663u,1.5 4459.538162662663u,0 4460.514702702702u,0 4460.515702702703u,1.5 4462.469782782783u,1.5 4462.470782782783u,0 4463.447322822823u,0 4463.448322822823u,1.5 4465.402402902902u,1.5 4465.403402902903u,0 4466.379942942943u,0 4466.380942942943u,1.5 4467.357482982983u,1.5 4467.358482982983u,0 4468.335023023023u,0 4468.336023023023u,1.5 4469.312563063063u,1.5 4469.313563063063u,0 4470.290103103103u,0 4470.2911031031035u,1.5 4471.267643143143u,1.5 4471.268643143143u,0 4472.245183183183u,0 4472.246183183183u,1.5 4473.222723223223u,1.5 4473.223723223223u,0 4476.155343343343u,0 4476.156343343343u,1.5 4478.1104234234235u,1.5 4478.111423423424u,0 4479.087963463464u,0 4479.088963463464u,1.5 4480.065503503503u,1.5 4480.066503503504u,0 4488.863363863864u,0 4488.864363863864u,1.5 4495.706144144144u,1.5 4495.707144144144u,0 4496.683684184184u,0 4496.684684184184u,1.5 4497.661224224224u,1.5 4497.662224224224u,0 4502.5489244244245u,0 4502.549924424425u,1.5 4503.526464464465u,1.5 4503.527464464465u,0 4504.504004504504u,0 4504.5050045045045u,1.5 4506.459084584585u,1.5 4506.460084584585u,0 4516.234484984985u,0 4516.235484984985u,1.5 4517.212025025025u,1.5 4517.213025025025u,0 4519.167105105105u,0 4519.1681051051055u,1.5 4520.144645145145u,1.5 4520.145645145145u,0 4521.122185185185u,0 4521.123185185185u,1.5 4523.077265265266u,1.5 4523.078265265266u,0 4524.054805305305u,0 4524.0558053053055u,1.5 4525.032345345345u,1.5 4525.033345345345u,0 4526.009885385385u,0 4526.010885385385u,1.5 4526.9874254254255u,1.5 4526.988425425426u,0 4528.942505505505u,0 4528.9435055055055u,1.5 4530.897585585586u,1.5 4530.898585585586u,0 4532.852665665666u,0 4532.853665665666u,1.5 4534.807745745745u,1.5 4534.808745745745u,0 4535.785285785786u,0 4535.786285785786u,1.5 4546.538226226226u,1.5 4546.539226226226u,0 4547.515766266267u,0 4547.516766266267u,1.5 4549.470846346346u,1.5 4549.471846346346u,0 4551.4259264264265u,0 4551.426926426427u,1.5 4552.403466466467u,1.5 4552.404466466467u,0 4556.3136266266265u,0 4556.314626626627u,1.5 4557.291166666667u,1.5 4557.292166666667u,0 4565.111486986987u,0 4565.112486986987u,1.5 4566.0890270270265u,1.5 4566.090027027027u,0 4567.066567067067u,0 4567.067567067067u,1.5 4571.954267267268u,1.5 4571.955267267268u,0 4572.931807307307u,0 4572.9328073073075u,1.5 4575.8644274274275u,1.5 4575.865427427428u,0 4576.841967467468u,0 4576.842967467468u,1.5 4577.819507507507u,1.5 4577.8205075075075u,0 4578.797047547547u,0 4578.798047547547u,1.5 4579.774587587588u,1.5 4579.775587587588u,0 4584.662287787788u,0 4584.663287787788u,1.5 4585.6398278278275u,1.5 4585.640827827828u,0 4586.617367867868u,0 4586.618367867868u,1.5 4597.370308308308u,1.5 4597.3713083083085u,0 4598.347848348348u,0 4598.348848348348u,1.5 4599.325388388388u,1.5 4599.326388388388u,0 4601.280468468469u,0 4601.281468468469u,1.5 4602.258008508508u,1.5 4602.2590085085085u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4609.100788788789u,1.5 4609.101788788789u,0 4610.0783288288285u,0 4610.079328828829u,1.5 4613.988488988989u,1.5 4613.989488988989u,0 4614.9660290290285u,0 4614.967029029029u,1.5 4615.943569069069u,1.5 4615.944569069069u,0 4616.921109109109u,0 4616.922109109109u,1.5 4617.898649149149u,1.5 4617.899649149149u,0 4620.83126926927u,0 4620.83226926927u,1.5 4623.763889389389u,1.5 4623.764889389389u,0 4624.741429429429u,0 4624.74242942943u,1.5 4627.674049549549u,1.5 4627.675049549549u,0 4630.60666966967u,0 4630.60766966967u,1.5 4631.584209709709u,1.5 4631.5852097097095u,0 4635.49436986987u,0 4635.49536986987u,1.5 4636.471909909909u,1.5 4636.4729099099095u,0 4637.44944994995u,0 4637.45044994995u,1.5 4641.35961011011u,1.5 4641.36061011011u,0 4642.33715015015u,0 4642.33815015015u,1.5 4643.31469019019u,1.5 4643.31569019019u,0 4644.2922302302295u,0 4644.29323023023u,1.5 4645.269770270271u,1.5 4645.270770270271u,0 4648.20239039039u,0 4648.20339039039u,1.5 4649.17993043043u,1.5 4649.180930430431u,0 4651.13501051051u,0 4651.1360105105105u,1.5 4656.02271071071u,1.5 4656.0237107107105u,0 4657.977790790791u,0 4657.978790790791u,1.5 4658.9553308308305u,1.5 4658.956330830831u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4667.753191191191u,1.5 4667.754191191191u,0 4675.573511511511u,0 4675.574511511511u,1.5 4680.461211711711u,1.5 4680.4622117117115u,0 4682.416291791792u,0 4682.417291791792u,1.5 4683.393831831831u,1.5 4683.394831831832u,0 4686.326451951952u,0 4686.327451951952u,1.5 4689.259072072072u,1.5 4689.260072072072u,0 4690.236612112112u,0 4690.237612112112u,1.5 4691.214152152152u,1.5 4691.215152152152u,0 4693.1692322322315u,0 4693.170232232232u,1.5 4694.146772272273u,1.5 4694.147772272273u,0 4696.101852352352u,0 4696.102852352352u,1.5 4698.056932432432u,1.5 4698.057932432433u,0 4699.034472472473u,0 4699.035472472473u,1.5 4700.012012512512u,1.5 4700.013012512512u,0 4703.922172672673u,0 4703.923172672673u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4712.720033033032u,1.5 4712.721033033033u,0 4715.652653153153u,0 4715.653653153153u,1.5 4717.6077332332325u,1.5 4717.608733233233u,0 4718.585273273274u,0 4718.586273273274u,1.5 4719.562813313313u,1.5 4719.563813313313u,0 4720.540353353353u,0 4720.541353353353u,1.5 4723.472973473474u,1.5 4723.473973473474u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4731.293293793794u,1.5 4731.294293793794u,0 4732.270833833833u,0 4732.271833833834u,1.5 4735.203453953954u,1.5 4735.204453953954u,0 4739.113614114114u,0 4739.114614114114u,1.5 4740.091154154154u,1.5 4740.092154154154u,0 4741.068694194194u,0 4741.069694194194u,1.5 4742.046234234233u,1.5 4742.047234234234u,0 4743.023774274275u,0 4743.024774274275u,1.5 4744.001314314314u,1.5 4744.002314314314u,0 4744.978854354354u,0 4744.979854354354u,1.5 4745.956394394394u,1.5 4745.957394394394u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4754.7542547547555u,1.5 4754.755254754756u,0 4755.731794794795u,0 4755.732794794795u,1.5 4756.709334834834u,1.5 4756.710334834835u,0 4759.6419549549555u,0 4759.642954954956u,1.5 4760.619494994995u,1.5 4760.620494994995u,0 4761.597035035034u,0 4761.598035035035u,1.5 4763.552115115115u,1.5 4763.553115115115u,0 4764.5296551551555u,0 4764.530655155156u,1.5 4765.507195195195u,1.5 4765.508195195195u,0 4767.462275275276u,0 4767.463275275276u,1.5 4769.4173553553555u,1.5 4769.418355355356u,0 4771.372435435435u,0 4771.373435435436u,1.5 4777.237675675676u,1.5 4777.238675675676u,0 4782.125375875876u,0 4782.126375875876u,1.5 4783.102915915916u,1.5 4783.103915915916u,0 4784.0804559559565u,0 4784.081455955957u,1.5 4787.990616116116u,1.5 4787.991616116116u,0 4793.8558563563565u,0 4793.856856356357u,1.5 4796.788476476477u,1.5 4796.789476476477u,0 4797.766016516516u,0 4797.767016516516u,1.5 4799.721096596597u,1.5 4799.722096596597u,0 4802.653716716716u,0 4802.654716716716u,1.5 4803.6312567567575u,1.5 4803.632256756758u,0 4807.541416916917u,0 4807.542416916917u,1.5 4809.496496996997u,1.5 4809.497496996997u,0 4815.361737237236u,0 4815.362737237237u,1.5 4819.271897397397u,1.5 4819.272897397397u,0 4820.249437437437u,0 4820.2504374374375u,1.5 4822.204517517517u,1.5 4822.205517517517u,0 4824.159597597598u,0 4824.160597597598u,1.5 4826.114677677678u,1.5 4826.115677677678u,0 4828.069757757758u,0 4828.070757757759u,1.5 4831.002377877878u,1.5 4831.003377877878u,0 4831.979917917918u,0 4831.980917917918u,1.5 4832.9574579579585u,1.5 4832.958457957959u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4840.777778278279u,1.5 4840.778778278279u,0 4842.7328583583585u,0 4842.733858358359u,1.5 4844.687938438438u,1.5 4844.6889384384385u,0 4848.598098598599u,0 4848.599098598599u,1.5 4849.575638638638u,1.5 4849.5766386386385u,0 4852.508258758759u,0 4852.50925875876u,1.5 4854.463338838838u,1.5 4854.464338838839u,0 4855.440878878879u,0 4855.441878878879u,1.5 4857.395958958959u,1.5 4857.39695895896u,0 4863.261199199199u,0 4863.262199199199u,1.5 4864.238739239238u,1.5 4864.239739239239u,0 4866.193819319319u,0 4866.194819319319u,1.5 4869.126439439439u,1.5 4869.1274394394395u,0 4870.10397947948u,0 4870.10497947948u,1.5 4871.081519519519u,1.5 4871.082519519519u,0 4872.0590595595595u,0 4872.06005955956u,1.5 4874.014139639639u,1.5 4874.0151396396395u,0 4875.969219719719u,0 4875.970219719719u,1.5 4876.94675975976u,1.5 4876.947759759761u,0 4877.9242997998u,0 4877.9252997998u,1.5 4878.901839839839u,1.5 4878.9028398398395u,0 4879.87937987988u,0 4879.88037987988u,1.5 4880.85691991992u,1.5 4880.85791991992u,0 4881.83445995996u,0 4881.835459959961u,1.5 4883.789540040039u,1.5 4883.79054004004u,0 4884.76708008008u,0 4884.76808008008u,1.5 4886.7221601601605u,1.5 4886.723160160161u,0 4888.677240240239u,0 4888.67824024024u,1.5 4889.654780280281u,1.5 4889.655780280281u,0 4891.6098603603605u,0 4891.610860360361u,1.5 4892.5874004004u,1.5 4892.5884004004u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4894.542480480481u,1.5 4894.543480480481u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4898.45264064064u,1.5 4898.4536406406405u,0 4899.430180680681u,0 4899.431180680681u,1.5 4900.40772072072u,1.5 4900.40872072072u,0 4901.385260760761u,0 4901.386260760762u,1.5 4903.34034084084u,1.5 4903.3413408408405u,0 4904.317880880881u,0 4904.318880880881u,1.5 4905.295420920921u,1.5 4905.296420920921u,0 4912.138201201201u,0 4912.139201201201u,1.5 4913.11574124124u,1.5 4913.116741241241u,0 4914.093281281282u,0 4914.094281281282u,1.5 4915.070821321321u,1.5 4915.071821321321u,0 4918.003441441441u,0 4918.0044414414415u,1.5 4919.958521521521u,1.5 4919.959521521521u,0 4920.9360615615615u,0 4920.937061561562u,1.5 4921.913601601602u,1.5 4921.914601601602u,0 4922.891141641641u,0 4922.8921416416415u,1.5 4923.868681681682u,1.5 4923.869681681682u,0 4925.823761761762u,0 4925.824761761763u,1.5 4926.801301801802u,1.5 4926.802301801802u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4938.531782282283u,0 4938.532782282283u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 4941.464402402402u,0 4941.465402402402u,1.5 4945.3745625625625u,1.5 4945.375562562563u,0 4946.352102602603u,0 4946.353102602603u,1.5 4947.329642642642u,1.5 4947.3306426426425u,0 4948.307182682683u,0 4948.308182682683u,1.5 4949.284722722722u,1.5 4949.285722722722u,0 4950.262262762763u,0 4950.263262762764u,1.5 4953.194882882883u,1.5 4953.195882882883u,0 4954.172422922923u,0 4954.173422922923u,1.5 4955.149962962963u,1.5 4955.150962962964u,0 4956.127503003003u,0 4956.128503003003u,1.5 4957.105043043042u,1.5 4957.1060430430425u,0 4965.902903403403u,0 4965.903903403403u,1.5 4966.880443443443u,1.5 4966.8814434434435u,0 4968.835523523523u,0 4968.836523523523u,1.5 4970.790603603604u,1.5 4970.791603603604u,0 4971.768143643643u,0 4971.7691436436435u,1.5 4972.745683683684u,1.5 4972.746683683684u,0 4973.723223723723u,0 4973.724223723723u,1.5 4974.700763763764u,1.5 4974.701763763765u,0 4975.678303803804u,0 4975.679303803804u,1.5 4976.655843843843u,1.5 4976.6568438438435u,0 4977.633383883884u,0 4977.634383883884u,1.5 4979.588463963964u,1.5 4979.589463963965u,0 4980.566004004004u,0 4980.567004004004u,1.5 4981.543544044043u,1.5 4981.5445440440435u,0 4982.521084084084u,0 4982.522084084084u,1.5 4983.498624124124u,1.5 4983.499624124124u,0 4984.476164164164u,0 4984.477164164165u,1.5 4986.431244244243u,1.5 4986.4322442442435u,0 4987.408784284285u,0 4987.409784284285u,1.5 4988.386324324324u,1.5 4988.387324324324u,0 4991.318944444444u,0 4991.319944444444u,1.5 4992.296484484485u,1.5 4992.297484484485u,0 4993.274024524524u,0 4993.275024524524u,1.5 4994.251564564564u,1.5 4994.252564564565u,0 4995.229104604605u,0 4995.230104604605u,1.5 4996.206644644644u,1.5 4996.2076446446445u,0 4998.161724724724u,0 4998.162724724724u,1.5 5007.937125125125u,1.5 5007.938125125125u,0 5009.892205205205u,0 5009.893205205205u,1.5 5014.779905405405u,1.5 5014.780905405405u,0 5015.757445445445u,0 5015.758445445445u,1.5 5016.734985485486u,1.5 5016.735985485486u,0 5017.712525525525u,0 5017.713525525525u,1.5 5021.622685685686u,1.5 5021.623685685686u,0 5022.600225725725u,0 5022.601225725725u,1.5 5024.555305805806u,1.5 5024.556305805806u,0 5025.532845845845u,0 5025.5338458458455u,1.5 5027.487925925926u,1.5 5027.488925925926u,0 5028.465465965966u,0 5028.466465965967u,1.5 5029.443006006006u,1.5 5029.444006006006u,0 5030.420546046045u,0 5030.4215460460455u,1.5 5031.398086086087u,1.5 5031.399086086087u,0 5033.353166166166u,0 5033.354166166167u,1.5 5035.308246246245u,1.5 5035.3092462462455u,0 5039.218406406406u,0 5039.219406406406u,1.5 5040.195946446446u,1.5 5040.196946446446u,0 5043.128566566566u,0 5043.129566566567u,1.5 5044.106106606607u,1.5 5044.107106606607u,0 5046.061186686687u,0 5046.062186686687u,1.5 5047.038726726726u,1.5 5047.039726726726u,0 5049.971346846846u,0 5049.972346846846u,1.5 5050.948886886887u,1.5 5050.949886886887u,0 5052.903966966967u,0 5052.904966966968u,1.5 5057.791667167167u,1.5 5057.792667167168u,0 5058.769207207207u,0 5058.770207207207u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5064.634447447447u,1.5 5064.635447447447u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5068.544607607608u,0 5068.545607607608u,1.5 5069.522147647647u,1.5 5069.523147647647u,0 5076.364927927928u,0 5076.365927927928u,1.5 5078.320008008008u,1.5 5078.321008008008u,0 5079.297548048047u,0 5079.298548048047u,1.5 5083.207708208208u,1.5 5083.208708208208u,0 5084.185248248248u,0 5084.186248248248u,1.5 5086.140328328328u,1.5 5086.141328328328u,0 5087.117868368368u,0 5087.118868368369u,1.5 5088.095408408408u,1.5 5088.096408408408u,0 5090.050488488489u,0 5090.051488488489u,1.5 5093.960648648648u,1.5 5093.961648648648u,0 5096.893268768769u,0 5096.8942687687695u,1.5 5097.870808808809u,1.5 5097.871808808809u,0 5098.848348848848u,0 5098.849348848848u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5112.533909409409u,0 5112.534909409409u,1.5 5113.511449449449u,1.5 5113.512449449449u,0 5114.4889894894895u,0 5114.48998948949u,1.5 5115.466529529529u,1.5 5115.467529529529u,0 5116.444069569569u,0 5116.44506956957u,1.5 5120.354229729729u,1.5 5120.355229729729u,0 5121.33176976977u,0 5121.3327697697705u,1.5 5123.286849849849u,1.5 5123.287849849849u,0 5124.26438988989u,0 5124.26538988989u,1.5 5125.24192992993u,1.5 5125.24292992993u,0 5128.174550050049u,0 5128.175550050049u,1.5 5129.1520900900905u,1.5 5129.153090090091u,0 5130.12963013013u,0 5130.13063013013u,1.5 5131.10717017017u,1.5 5131.1081701701705u,0 5132.08471021021u,0 5132.08571021021u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5135.99487037037u,0 5135.9958703703705u,1.5 5136.97241041041u,1.5 5136.97341041041u,0 5142.83765065065u,0 5142.83865065065u,1.5 5143.8151906906905u,1.5 5143.816190690691u,0 5144.79273073073u,0 5144.79373073073u,1.5 5149.680430930931u,1.5 5149.681430930931u,0 5150.657970970971u,0 5150.6589709709715u,1.5 5152.61305105105u,1.5 5152.61405105105u,0 5153.5905910910915u,0 5153.591591091092u,1.5 5156.523211211211u,1.5 5156.524211211211u,0 5157.500751251251u,0 5157.501751251251u,1.5 5158.4782912912915u,1.5 5158.479291291292u,0 5159.455831331331u,0 5159.456831331331u,1.5 5160.433371371371u,1.5 5160.4343713713715u,0 5161.410911411411u,0 5161.411911411411u,1.5 5162.388451451451u,1.5 5162.389451451451u,0 5168.2536916916915u,0 5168.254691691692u,1.5 5170.208771771772u,1.5 5170.2097717717725u,0 5172.163851851851u,0 5172.164851851851u,1.5 5174.118931931932u,1.5 5174.119931931932u,0 5176.074012012012u,0 5176.075012012012u,1.5 5177.051552052051u,1.5 5177.052552052051u,0 5181.939252252252u,0 5181.940252252252u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5190.737112612613u,0 5190.738112612613u,1.5 5193.669732732732u,1.5 5193.670732732732u,0 5195.624812812813u,0 5195.625812812813u,1.5 5198.557432932933u,1.5 5198.558432932933u,0 5199.534972972973u,0 5199.5359729729735u,1.5 5200.512513013013u,1.5 5200.513513013013u,0 5201.490053053052u,0 5201.491053053052u,1.5 5202.4675930930935u,1.5 5202.468593093094u,0 5203.445133133133u,0 5203.446133133133u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5213.220533533533u,0 5213.221533533533u,1.5 5218.108233733733u,1.5 5218.109233733733u,0 5220.063313813814u,0 5220.064313813814u,1.5 5221.040853853853u,1.5 5221.041853853853u,0 5222.995933933934u,0 5222.996933933934u,1.5 5223.973473973974u,1.5 5223.974473973974u,0 5225.928554054053u,0 5225.929554054053u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5232.771334334334u,1.5 5232.772334334334u,0 5235.703954454454u,0 5235.704954454454u,1.5 5237.659034534534u,1.5 5237.660034534534u,0 5238.636574574574u,0 5238.6375745745745u,1.5 5240.591654654654u,1.5 5240.592654654654u,0 5244.501814814815u,0 5244.502814814815u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5254.277215215215u,0 5254.278215215215u,1.5 5255.254755255255u,1.5 5255.255755255255u,0 5256.232295295295u,0 5256.233295295296u,1.5 5258.187375375375u,1.5 5258.1883753753755u,0 5261.1199954954955u,0 5261.120995495496u,1.5 5262.097535535535u,1.5 5262.098535535535u,0 5266.0076956956955u,0 5266.008695695696u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5275.783096096096u,0 5275.784096096097u,1.5 5276.760636136136u,1.5 5276.761636136136u,0 5277.738176176176u,0 5277.739176176176u,1.5 5280.670796296296u,1.5 5280.671796296297u,0 5281.648336336336u,0 5281.649336336336u,1.5 5282.625876376376u,1.5 5282.6268763763765u,0 5283.603416416417u,0 5283.604416416417u,1.5 5285.558496496496u,1.5 5285.559496496497u,0 5287.513576576576u,0 5287.5145765765765u,1.5 5288.491116616617u,1.5 5288.492116616617u,0 5290.4461966966965u,0 5290.447196696697u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5294.356356856857u,0 5294.357356856857u,1.5 5295.3338968968965u,1.5 5295.334896896897u,0 5296.311436936937u,0 5296.312436936937u,1.5 5297.288976976977u,1.5 5297.289976976977u,0 5300.221597097097u,0 5300.222597097098u,1.5 5302.176677177177u,1.5 5302.177677177177u,0 5303.154217217217u,0 5303.155217217217u,1.5 5304.131757257258u,1.5 5304.132757257258u,0 5305.109297297297u,0 5305.110297297298u,1.5 5306.086837337337u,1.5 5306.087837337337u,0 5307.064377377377u,0 5307.065377377377u,1.5 5308.041917417418u,1.5 5308.042917417418u,0 5309.019457457458u,0 5309.020457457458u,1.5 5312.929617617618u,1.5 5312.930617617618u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5320.749937937938u,0 5320.750937937938u,1.5 5322.705018018018u,1.5 5322.706018018018u,0 5323.682558058058u,0 5323.683558058058u,1.5 5326.615178178178u,1.5 5326.616178178178u,0 5327.592718218218u,0 5327.593718218218u,1.5 5329.547798298298u,1.5 5329.548798298299u,0 5330.525338338338u,0 5330.526338338338u,1.5 5331.502878378378u,1.5 5331.503878378378u,0 5332.480418418419u,0 5332.481418418419u,1.5 5334.435498498498u,1.5 5334.436498498499u,0 5335.413038538538u,0 5335.414038538538u,1.5 5337.368118618619u,1.5 5337.369118618619u,0 5338.345658658659u,0 5338.346658658659u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5344.210898898898u,0 5344.211898898899u,1.5 5353.00875925926u,1.5 5353.00975925926u,0 5354.963839339339u,0 5354.964839339339u,1.5 5356.91891941942u,1.5 5356.91991941942u,0 5357.89645945946u,0 5357.89745945946u,1.5 5361.80661961962u,1.5 5361.80761961962u,0 5363.761699699699u,0 5363.7626996997u,1.5 5364.739239739739u,1.5 5364.740239739739u,0 5366.69431981982u,0 5366.69531981982u,1.5 5368.649399899899u,1.5 5368.6503998999u,0 5371.58202002002u,0 5371.58302002002u,1.5 5374.51464014014u,1.5 5374.51564014014u,0 5375.49218018018u,0 5375.49318018018u,1.5 5376.46972022022u,1.5 5376.47072022022u,0 5377.447260260261u,0 5377.448260260261u,1.5 5378.4248003003u,1.5 5378.425800300301u,0 5386.245120620621u,0 5386.246120620621u,1.5 5394.065440940941u,1.5 5394.066440940941u,0 5395.042980980981u,0 5395.043980980981u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5396.998061061061u,0 5396.999061061061u,1.5 5397.975601101101u,1.5 5397.976601101102u,0 5398.953141141141u,0 5398.954141141141u,1.5 5399.930681181181u,1.5 5399.931681181181u,0 5400.908221221221u,0 5400.909221221221u,1.5 5401.885761261262u,1.5 5401.886761261262u,0 5402.863301301301u,0 5402.864301301302u,1.5 5406.773461461462u,1.5 5406.774461461462u,0 5408.728541541541u,0 5408.729541541541u,1.5 5409.706081581581u,1.5 5409.707081581581u,0 5411.661161661662u,0 5411.662161661662u,1.5 5413.616241741741u,1.5 5413.617241741741u,0 5421.436562062062u,0 5421.437562062062u,1.5 5422.414102102102u,1.5 5422.4151021021025u,0 5424.369182182182u,0 5424.370182182182u,1.5 5425.346722222222u,1.5 5425.347722222222u,0 5426.324262262263u,0 5426.325262262263u,1.5 5429.256882382382u,1.5 5429.257882382382u,0 5431.211962462463u,0 5431.212962462463u,1.5 5432.189502502502u,1.5 5432.190502502503u,0 5433.167042542542u,0 5433.168042542542u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5438.054742742742u,0 5438.055742742742u,1.5 5439.032282782783u,1.5 5439.033282782783u,0 5440.009822822823u,0 5440.010822822823u,1.5 5440.987362862863u,1.5 5440.988362862863u,0 5443.919982982983u,0 5443.920982982983u,1.5 5445.875063063063u,1.5 5445.876063063063u,0 5446.852603103103u,0 5446.8536031031035u,1.5 5447.830143143143u,1.5 5447.831143143143u,0 5448.807683183183u,0 5448.808683183183u,1.5 5450.762763263264u,1.5 5450.763763263264u,0 5451.740303303303u,0 5451.7413033033035u,1.5 5457.605543543543u,1.5 5457.606543543543u,0 5458.583083583583u,0 5458.584083583583u,1.5 5461.515703703703u,1.5 5461.516703703704u,0 5462.493243743743u,0 5462.494243743743u,1.5 5464.448323823824u,1.5 5464.449323823824u,0 5465.425863863864u,0 5465.426863863864u,1.5 5470.313564064064u,1.5 5470.314564064064u,0 5471.291104104104u,0 5471.2921041041045u,1.5 5473.246184184184u,1.5 5473.247184184184u,0 5474.223724224224u,0 5474.224724224224u,1.5 5475.201264264265u,1.5 5475.202264264265u,0 5478.133884384384u,0 5478.134884384384u,1.5 5479.1114244244245u,1.5 5479.112424424425u,0 5480.088964464465u,0 5480.089964464465u,1.5 5482.044044544544u,1.5 5482.045044544544u,0 5483.021584584585u,0 5483.022584584585u,1.5 5485.954204704704u,1.5 5485.955204704705u,0 5486.931744744744u,0 5486.932744744744u,1.5 5487.909284784785u,1.5 5487.910284784785u,0 5488.8868248248245u,0 5488.887824824825u,1.5 5489.864364864865u,1.5 5489.865364864865u,0 5490.841904904904u,0 5490.842904904905u,1.5 5491.819444944945u,1.5 5491.820444944945u,0 5492.796984984985u,0 5492.797984984985u,1.5 5494.752065065065u,1.5 5494.753065065065u,0 5495.729605105105u,0 5495.7306051051055u,1.5 5496.707145145145u,1.5 5496.708145145145u,0 5499.639765265266u,0 5499.640765265266u,1.5 5500.617305305305u,1.5 5500.6183053053055u,0 5503.5499254254255u,0 5503.550925425426u,1.5 5504.527465465466u,1.5 5504.528465465466u,0 5509.415165665666u,0 5509.416165665666u,1.5 5512.347785785786u,1.5 5512.348785785786u,0 5515.280405905905u,0 5515.281405905906u,1.5 5516.257945945946u,1.5 5516.258945945946u,0 5517.235485985986u,0 5517.236485985986u,1.5 5518.213026026026u,1.5 5518.214026026026u,0 5520.168106106106u,0 5520.1691061061065u,1.5 5521.145646146146u,1.5 5521.146646146146u,0 5524.078266266267u,0 5524.079266266267u,1.5 5525.055806306306u,1.5 5525.0568063063065u,0 5526.033346346346u,0 5526.034346346346u,1.5 5527.010886386386u,1.5 5527.011886386386u,0 5527.9884264264265u,0 5527.989426426427u,1.5 5529.943506506506u,1.5 5529.9445065065065u,0 5530.921046546546u,0 5530.922046546546u,1.5 5531.898586586587u,1.5 5531.899586586587u,0 5533.853666666667u,0 5533.854666666667u,1.5 5538.741366866867u,1.5 5538.742366866867u,0 5539.718906906906u,0 5539.7199069069065u,1.5 5540.696446946947u,1.5 5540.697446946947u,0 5541.673986986987u,0 5541.674986986987u,1.5 5542.6515270270265u,1.5 5542.652527027027u,0 5543.629067067067u,0 5543.630067067067u,1.5 5547.539227227227u,1.5 5547.540227227227u,0 5548.516767267268u,0 5548.517767267268u,1.5 5549.494307307307u,1.5 5549.4953073073075u,0 5550.471847347347u,0 5550.472847347347u,1.5 5552.4269274274275u,1.5 5552.427927427428u,0 5557.3146276276275u,0 5557.315627627628u,1.5 5560.247247747748u,1.5 5560.248247747748u,0 5562.2023278278275u,0 5562.203327827828u,1.5 5563.179867867868u,1.5 5563.180867867868u,0 5566.112487987988u,0 5566.113487987988u,1.5 5567.0900280280275u,1.5 5567.091028028028u,0 5568.067568068068u,0 5568.068568068068u,1.5 5570.022648148148u,1.5 5570.023648148148u,0 5571.000188188188u,0 5571.001188188188u,1.5 5572.955268268269u,1.5 5572.956268268269u,0 5573.932808308308u,0 5573.9338083083085u,1.5 5575.887888388388u,1.5 5575.888888388388u,0 5577.842968468469u,0 5577.843968468469u,1.5 5578.820508508508u,1.5 5578.8215085085085u,0 5579.798048548548u,0 5579.799048548548u,1.5 5580.775588588589u,1.5 5580.776588588589u,0 5584.685748748749u,0 5584.686748748749u,1.5 5585.663288788789u,1.5 5585.664288788789u,0 5586.6408288288285u,0 5586.641828828829u,1.5 5587.618368868869u,1.5 5587.619368868869u,0 5589.573448948949u,0 5589.574448948949u,1.5 5595.438689189189u,1.5 5595.439689189189u,0 5596.4162292292285u,0 5596.417229229229u,1.5 5597.39376926927u,1.5 5597.39476926927u,0 5600.326389389389u,0 5600.327389389389u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5605.21408958959u,0 5605.21508958959u,1.5 5608.146709709709u,1.5 5608.1477097097095u,0 5609.12424974975u,0 5609.12524974975u,1.5 5610.10178978979u,1.5 5610.10278978979u,0 5611.0793298298295u,0 5611.08032982983u,1.5 5613.034409909909u,1.5 5613.0354099099095u,0 5614.01194994995u,0 5614.01294994995u,1.5 5614.98948998999u,1.5 5614.99048998999u,0 5615.9670300300295u,0 5615.96803003003u,1.5 5616.94457007007u,1.5 5616.94557007007u,0 5620.8547302302295u,0 5620.85573023023u,1.5 5621.832270270271u,1.5 5621.833270270271u,0 5623.78735035035u,0 5623.78835035035u,1.5 5628.67505055055u,1.5 5628.67605055055u,0 5629.652590590591u,0 5629.653590590591u,1.5 5630.63013063063u,1.5 5630.631130630631u,0 5632.58521071071u,0 5632.5862107107105u,1.5 5634.540290790791u,1.5 5634.541290790791u,0 5636.495370870871u,0 5636.496370870871u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5638.450450950951u,0 5638.451450950951u,1.5 5641.383071071071u,1.5 5641.384071071071u,0 5642.360611111111u,0 5642.361611111111u,1.5 5644.315691191191u,1.5 5644.316691191191u,0 5648.225851351351u,0 5648.226851351351u,1.5 5649.203391391391u,1.5 5649.204391391391u,0 5650.180931431431u,0 5650.181931431432u,1.5 5651.158471471472u,1.5 5651.159471471472u,0 5652.136011511511u,0 5652.137011511511u,1.5 5653.113551551551u,1.5 5653.114551551551u,0 5655.068631631631u,0 5655.069631631632u,1.5 5657.023711711711u,1.5 5657.0247117117115u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5664.8440320320315u,1.5 5664.845032032032u,0 5665.821572072072u,0 5665.822572072072u,1.5 5666.799112112112u,1.5 5666.800112112112u,0 5667.776652152152u,0 5667.777652152152u,1.5 5669.7317322322315u,1.5 5669.732732232232u,0 5675.596972472473u,0 5675.597972472473u,1.5 5676.574512512512u,1.5 5676.575512512512u,0 5678.529592592593u,0 5678.530592592593u,1.5 5679.507132632632u,1.5 5679.508132632633u,0 5680.484672672673u,0 5680.485672672673u,1.5 5683.417292792793u,1.5 5683.418292792793u,0 5684.394832832832u,0 5684.395832832833u,1.5 5688.304992992993u,1.5 5688.305992992993u,0 5689.282533033032u,0 5689.283533033033u,1.5 5690.260073073073u,1.5 5690.261073073073u,0 5691.237613113113u,0 5691.238613113113u,1.5 5692.215153153153u,1.5 5692.216153153153u,0 5695.147773273274u,0 5695.148773273274u,1.5 5696.125313313313u,1.5 5696.126313313313u,0 5699.057933433433u,0 5699.058933433434u,1.5 5700.035473473474u,1.5 5700.036473473474u,0 5701.013013513513u,0 5701.014013513513u,1.5 5702.968093593594u,1.5 5702.969093593594u,0 5703.945633633633u,0 5703.946633633634u,1.5 5704.923173673674u,1.5 5704.924173673674u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5711.765953953954u,1.5 5711.766953953954u,0 5713.721034034033u,0 5713.722034034034u,1.5 5716.653654154154u,1.5 5716.654654154154u,0 5718.608734234233u,0 5718.609734234234u,1.5 5722.518894394394u,1.5 5722.519894394394u,0 5723.496434434434u,0 5723.497434434435u,1.5 5725.451514514514u,1.5 5725.452514514514u,0 5726.429054554554u,0 5726.430054554554u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5734.249374874875u,1.5 5734.250374874875u,0 5740.114615115115u,0 5740.115615115115u,1.5 5744.024775275276u,1.5 5744.025775275276u,0 5745.002315315315u,0 5745.003315315315u,1.5 5746.957395395395u,1.5 5746.958395395395u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 5755.7552557557565u,1.5 5755.756255755757u,0 5757.710335835835u,0 5757.711335835836u,1.5 5759.665415915916u,1.5 5759.666415915916u,0 5760.6429559559565u,0 5760.643955955957u,1.5 5761.620495995996u,1.5 5761.621495995996u,0 5762.598036036035u,0 5762.599036036036u,1.5 5764.553116116116u,1.5 5764.554116116116u,0 5766.508196196196u,0 5766.509196196196u,1.5 5767.485736236235u,1.5 5767.486736236236u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5772.373436436436u,0 5772.374436436437u,1.5 5775.3060565565565u,1.5 5775.307056556557u,0 5776.283596596597u,0 5776.284596596597u,1.5 5777.261136636636u,1.5 5777.262136636637u,0 5778.238676676677u,0 5778.239676676677u,1.5 5779.216216716716u,1.5 5779.217216716716u,0 5780.1937567567575u,0 5780.194756756758u,1.5 5782.148836836836u,1.5 5782.149836836837u,0 5783.126376876877u,0 5783.127376876877u,1.5 5785.0814569569575u,1.5 5785.082456956958u,0 5786.058996996997u,0 5786.059996996997u,1.5 5787.036537037036u,1.5 5787.037537037037u,0 5788.014077077077u,0 5788.015077077077u,1.5 5792.901777277278u,1.5 5792.902777277278u,0 5793.879317317317u,0 5793.880317317317u,1.5 5794.8568573573575u,1.5 5794.857857357358u,0 5795.834397397397u,0 5795.835397397397u,1.5 5798.767017517517u,1.5 5798.768017517517u,0 5799.7445575575575u,0 5799.745557557558u,1.5 5801.699637637637u,1.5 5801.700637637638u,0 5802.677177677678u,0 5802.678177677678u,1.5 5809.5199579579585u,1.5 5809.520957957959u,0 5813.430118118118u,0 5813.431118118118u,1.5 5815.385198198198u,1.5 5815.386198198198u,0 5817.340278278279u,0 5817.341278278279u,1.5 5821.250438438438u,1.5 5821.2514384384385u,0 5822.227978478479u,0 5822.228978478479u,1.5 5823.205518518518u,1.5 5823.206518518518u,0 5825.160598598599u,0 5825.161598598599u,1.5 5827.115678678679u,1.5 5827.116678678679u,0 5829.070758758759u,0 5829.07175875876u,1.5 5830.048298798799u,1.5 5830.049298798799u,0 5831.025838838838u,0 5831.026838838839u,1.5 5833.958458958959u,1.5 5833.95945895896u,0 5837.868619119119u,0 5837.869619119119u,1.5 5838.8461591591595u,1.5 5838.84715915916u,0 5840.801239239238u,0 5840.802239239239u,1.5 5842.756319319319u,1.5 5842.757319319319u,0 5843.7338593593595u,0 5843.73485935936u,1.5 5845.688939439439u,1.5 5845.6899394394395u,0 5849.5990995996u,0 5849.6000995996u,1.5 5851.55417967968u,1.5 5851.55517967968u,0 5852.531719719719u,0 5852.532719719719u,1.5 5856.44187987988u,1.5 5856.44287987988u,0 5858.39695995996u,0 5858.397959959961u,1.5 5860.352040040039u,1.5 5860.35304004004u,0 5862.30712012012u,0 5862.30812012012u,1.5 5871.104980480481u,1.5 5871.105980480481u,0 5872.08252052052u,0 5872.08352052052u,1.5 5873.0600605605605u,1.5 5873.061060560561u,0 5876.97022072072u,0 5876.97122072072u,1.5 5877.947760760761u,1.5 5877.948760760762u,0 5878.925300800801u,0 5878.926300800801u,1.5 5880.880380880881u,1.5 5880.881380880881u,0 5882.835460960961u,0 5882.836460960962u,1.5 5883.813001001001u,1.5 5883.814001001001u,0 5884.79054104104u,0 5884.791541041041u,1.5 5885.768081081081u,1.5 5885.769081081081u,0 5886.745621121121u,0 5886.746621121121u,1.5 5889.67824124124u,1.5 5889.679241241241u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5899.453641641641u,1.5 5899.4546416416415u,0 5901.408721721721u,0 5901.409721721721u,1.5 5903.363801801802u,1.5 5903.364801801802u,0 5906.296421921922u,0 5906.297421921922u,1.5 5907.273961961962u,1.5 5907.274961961963u,0 5908.251502002002u,0 5908.252502002002u,1.5 5911.184122122122u,1.5 5911.185122122122u,0 5912.161662162162u,0 5912.162662162163u,1.5 5920.959522522522u,1.5 5920.960522522522u,0 5921.9370625625625u,0 5921.938062562563u,1.5 5922.914602602603u,1.5 5922.915602602603u,0 5923.892142642642u,0 5923.8931426426425u,1.5 5924.869682682683u,1.5 5924.870682682683u,0 5925.847222722722u,0 5925.848222722722u,1.5 5926.824762762763u,1.5 5926.825762762764u,0 5931.712462962963u,0 5931.713462962964u,1.5 5933.667543043042u,1.5 5933.6685430430425u,0 5935.622623123123u,0 5935.623623123123u,1.5 5936.600163163163u,1.5 5936.601163163164u,0 5938.555243243242u,0 5938.5562432432425u,1.5 5946.375563563563u,1.5 5946.376563563564u,0 5947.353103603604u,0 5947.354103603604u,1.5 5948.330643643643u,1.5 5948.3316436436435u,0 5949.308183683684u,0 5949.309183683684u,1.5 5950.285723723723u,1.5 5950.286723723723u,0 5951.263263763764u,0 5951.264263763765u,1.5 5952.240803803804u,1.5 5952.241803803804u,0 5953.218343843843u,0 5953.2193438438435u,1.5 5954.195883883884u,1.5 5954.196883883884u,0 5957.128504004004u,0 5957.129504004004u,1.5 5959.083584084084u,1.5 5959.084584084084u,0 5960.061124124124u,0 5960.062124124124u,1.5 5961.038664164164u,1.5 5961.039664164165u,0 5962.993744244243u,0 5962.9947442442435u,1.5 5964.948824324324u,1.5 5964.949824324324u,0 5968.858984484485u,0 5968.859984484485u,1.5 5970.814064564564u,1.5 5970.815064564565u,0 5971.791604604605u,0 5971.792604604605u,1.5 5972.769144644644u,1.5 5972.7701446446445u,0 5973.746684684685u,0 5973.747684684685u,1.5 5979.611924924925u,1.5 5979.612924924925u,0 5980.589464964965u,0 5980.590464964966u,1.5 5983.522085085086u,1.5 5983.523085085086u,0 5984.499625125125u,0 5984.500625125125u,1.5 5986.454705205205u,1.5 5986.455705205205u,0 5987.432245245244u,0 5987.4332452452445u,1.5 6006.005506006006u,1.5 6006.006506006006u,0 6006.983046046045u,0 6006.9840460460455u,1.5 6012.848286286287u,1.5 6012.849286286287u,0 6013.825826326326u,0 6013.826826326326u,1.5 6017.735986486487u,1.5 6017.736986486487u,0 6018.713526526526u,0 6018.714526526526u,1.5 6023.601226726726u,1.5 6023.602226726726u,0 6024.578766766767u,0 6024.5797667667675u,1.5 6028.488926926927u,1.5 6028.489926926927u,0 6029.466466966967u,0 6029.467466966968u,1.5 6030.444007007007u,1.5 6030.445007007007u,0 6032.3990870870875u,0 6032.400087087088u,1.5 6033.376627127127u,1.5 6033.377627127127u,0 6036.309247247247u,0 6036.310247247247u,1.5 6038.264327327327u,1.5 6038.265327327327u,0 6044.129567567567u,0 6044.130567567568u,1.5 6045.107107607608u,1.5 6045.108107607608u,0 6049.994807807808u,0 6049.995807807808u,1.5 6054.882508008008u,1.5 6054.883508008008u,0 6057.815128128128u,0 6057.816128128128u,1.5 6059.770208208208u,1.5 6059.771208208208u,0 6060.747748248248u,0 6060.748748248248u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6068.568068568568u,0 6068.569068568569u,1.5 6073.455768768769u,1.5 6073.4567687687695u,0 6074.433308808809u,0 6074.434308808809u,1.5 6075.410848848848u,1.5 6075.411848848848u,0 6076.388388888889u,0 6076.389388888889u,1.5 6077.365928928929u,1.5 6077.366928928929u,0 6078.343468968969u,0 6078.3444689689695u,1.5 6079.321009009009u,1.5 6079.322009009009u,0 6080.298549049048u,0 6080.299549049048u,1.5 6087.141329329329u,1.5 6087.142329329329u,0 6088.118869369369u,0 6088.11986936937u,1.5 6090.073949449449u,1.5 6090.074949449449u,0 6095.93918968969u,0 6095.94018968969u,1.5 6096.916729729729u,1.5 6096.917729729729u,0 6097.89426976977u,0 6097.8952697697705u,1.5 6100.82688988989u,1.5 6100.82788988989u,0 6102.78196996997u,0 6102.7829699699705u,1.5 6103.75951001001u,1.5 6103.76051001001u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6106.69213013013u,1.5 6106.69313013013u,0 6107.66967017017u,0 6107.6706701701705u,1.5 6108.64721021021u,1.5 6108.64821021021u,0 6113.53491041041u,0 6113.53591041041u,1.5 6117.44507057057u,1.5 6117.446070570571u,0 6130.1530910910915u,0 6130.154091091092u,1.5 6136.018331331331u,1.5 6136.019331331331u,0 6137.973411411411u,0 6137.974411411411u,1.5 6141.883571571571u,1.5 6141.8845715715715u,0 6143.838651651651u,0 6143.839651651651u,1.5 6147.748811811812u,1.5 6147.749811811812u,0 6148.726351851851u,0 6148.727351851851u,1.5 6153.614052052051u,1.5 6153.615052052051u,0 6155.569132132132u,0 6155.570132132132u,1.5 6156.546672172172u,1.5 6156.5476721721725u,0 6157.524212212212u,0 6157.525212212212u,1.5 6158.501752252252u,1.5 6158.502752252252u,0 6160.456832332332u,0 6160.457832332332u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6168.277152652652u,0 6168.278152652652u,1.5 6171.209772772773u,1.5 6171.210772772773u,0 6173.164852852852u,0 6173.165852852852u,1.5 6175.119932932933u,1.5 6175.120932932933u,0 6176.097472972973u,0 6176.0984729729735u,1.5 6177.075013013013u,1.5 6177.076013013013u,0 6178.052553053052u,0 6178.053553053052u,1.5 6179.0300930930935u,1.5 6179.031093093094u,0 6180.985173173173u,0 6180.9861731731735u,1.5 6181.962713213213u,1.5 6181.963713213213u,0 6182.940253253253u,0 6182.941253253253u,1.5 6184.895333333333u,1.5 6184.896333333333u,0 6185.872873373373u,0 6185.8738733733735u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6190.760573573573u,0 6190.7615735735735u,1.5 6191.738113613614u,1.5 6191.739113613614u,0 6192.715653653653u,0 6192.716653653653u,1.5 6197.603353853853u,1.5 6197.604353853853u,0 6200.535973973974u,0 6200.536973973974u,1.5 6202.491054054053u,1.5 6202.492054054053u,0 6203.468594094094u,0 6203.469594094095u,1.5 6208.3562942942945u,1.5 6208.357294294295u,0 6213.2439944944945u,0 6213.244994494495u,1.5 6215.199074574574u,1.5 6215.2000745745745u,0 6216.176614614615u,0 6216.177614614615u,1.5 6219.109234734734u,1.5 6219.110234734734u,0 6220.086774774775u,0 6220.087774774775u,1.5 6222.041854854854u,1.5 6222.042854854854u,0 6223.0193948948945u,0 6223.020394894895u,1.5 6223.996934934935u,1.5 6223.997934934935u,0 6224.974474974975u,0 6224.975474974975u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6231.817255255255u,0 6231.818255255255u,1.5 6233.772335335335u,1.5 6233.773335335335u,0 6235.727415415415u,0 6235.728415415415u,1.5 6238.660035535535u,1.5 6238.661035535535u,0 6244.525275775776u,0 6244.526275775776u,1.5 6245.502815815816u,1.5 6245.503815815816u,0 6246.480355855855u,0 6246.481355855855u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6254.300676176176u,1.5 6254.301676176176u,0 6258.210836336336u,0 6258.211836336336u,1.5 6260.165916416417u,1.5 6260.166916416417u,0 6261.143456456457u,0 6261.144456456457u,1.5 6262.120996496496u,1.5 6262.121996496497u,0 6265.053616616617u,0 6265.054616616617u,1.5 6266.031156656657u,1.5 6266.032156656657u,0 6267.0086966966965u,0 6267.009696696697u,1.5 6268.963776776777u,1.5 6268.964776776777u,0 6269.941316816817u,0 6269.942316816817u,1.5 6270.918856856857u,1.5 6270.919856856857u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6273.851476976977u,1.5 6273.852476976977u,0 6274.829017017017u,0 6274.830017017017u,1.5 6275.806557057057u,1.5 6275.807557057057u,0 6276.784097097097u,0 6276.785097097098u,1.5 6277.761637137137u,1.5 6277.762637137137u,0 6279.716717217217u,0 6279.717717217217u,1.5 6282.649337337337u,1.5 6282.650337337337u,0 6283.626877377377u,0 6283.627877377377u,1.5 6284.604417417418u,1.5 6284.605417417418u,0 6287.537037537537u,0 6287.538037537537u,1.5 6288.514577577577u,1.5 6288.5155775775775u,0 6296.3348978978975u,0 6296.335897897898u,1.5 6298.289977977978u,1.5 6298.290977977978u,0 6300.245058058058u,0 6300.246058058058u,1.5 6304.155218218218u,1.5 6304.156218218218u,0 6305.132758258259u,0 6305.133758258259u,1.5 6309.042918418419u,1.5 6309.043918418419u,0 6310.020458458459u,0 6310.021458458459u,1.5 6313.930618618619u,1.5 6313.931618618619u,0 6314.908158658659u,0 6314.909158658659u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6317.840778778779u,0 6317.841778778779u,1.5 6318.818318818819u,1.5 6318.819318818819u,0 6319.795858858859u,0 6319.796858858859u,1.5 6320.773398898898u,1.5 6320.774398898899u,0 6321.750938938939u,0 6321.751938938939u,1.5 6326.638639139139u,1.5 6326.639639139139u,0 6329.57125925926u,0 6329.57225925926u,1.5 6330.548799299299u,1.5 6330.5497992993u,0 6331.526339339339u,0 6331.527339339339u,1.5 6337.391579579579u,1.5 6337.392579579579u,0 6339.34665965966u,0 6339.34765965966u,1.5 6340.324199699699u,1.5 6340.3251996997u,0 6342.27927977978u,0 6342.28027977978u,1.5 6343.25681981982u,1.5 6343.25781981982u,0 6344.23435985986u,0 6344.23535985986u,1.5 6350.0996001001u,1.5 6350.100600100101u,0 6351.07714014014u,0 6351.07814014014u,1.5 6352.05468018018u,1.5 6352.05568018018u,0 6354.009760260261u,0 6354.010760260261u,1.5 6354.9873003003u,1.5 6354.988300300301u,0 6355.96484034034u,0 6355.96584034034u,1.5 6356.94238038038u,1.5 6356.94338038038u,0 6358.897460460461u,0 6358.898460460461u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6363.785160660661u,1.5 6363.786160660661u,0 6370.627940940941u,0 6370.628940940941u,1.5 6371.605480980981u,1.5 6371.606480980981u,0 6372.583021021021u,0 6372.584021021021u,1.5 6379.425801301301u,1.5 6379.426801301302u,0 6386.268581581581u,0 6386.269581581581u,1.5 6388.223661661662u,1.5 6388.224661661662u,0 6389.201201701701u,0 6389.202201701702u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6397.999062062062u,0 6398.000062062062u,1.5 6398.976602102102u,1.5 6398.9776021021025u,0 6400.931682182182u,0 6400.932682182182u,1.5 6401.909222222222u,1.5 6401.910222222222u,0 6404.841842342342u,0 6404.842842342342u,1.5 6406.7969224224225u,1.5 6406.797922422423u,0 6407.774462462463u,0 6407.775462462463u,1.5 6410.707082582582u,1.5 6410.708082582582u,0 6411.684622622623u,0 6411.685622622623u,1.5 6414.617242742742u,1.5 6414.618242742742u,0 6416.572322822823u,0 6416.573322822823u,1.5 6417.549862862863u,1.5 6417.550862862863u,0 6420.482482982983u,0 6420.483482982983u,1.5 6421.460023023023u,1.5 6421.461023023023u,0 6422.437563063063u,0 6422.438563063063u,1.5 6426.347723223223u,1.5 6426.348723223223u,0 6427.325263263264u,0 6427.326263263264u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6437.100663663664u,1.5 6437.101663663664u,0 6445.898524024024u,0 6445.899524024024u,1.5 6448.831144144144u,1.5 6448.832144144144u,0 6449.808684184184u,0 6449.809684184184u,1.5 6451.763764264265u,1.5 6451.764764264265u,0 6452.741304304304u,0 6452.7423043043045u,1.5 6454.696384384384u,1.5 6454.697384384384u,0 6456.651464464465u,0 6456.652464464465u,1.5 6463.494244744744u,1.5 6463.495244744744u,0 6464.471784784785u,0 6464.472784784785u,1.5 6465.4493248248245u,1.5 6465.450324824825u,0 6466.426864864865u,0 6466.427864864865u,1.5 6468.381944944945u,1.5 6468.382944944945u,0 6469.359484984985u,0 6469.360484984985u,1.5 6471.314565065065u,1.5 6471.315565065065u,0 6472.292105105105u,0 6472.2931051051055u,1.5 6474.247185185185u,1.5 6474.248185185185u,0 6476.202265265266u,0 6476.203265265266u,1.5 6477.179805305305u,1.5 6477.1808053053055u,0 6484.022585585586u,0 6484.023585585586u,1.5 6485.0001256256255u,1.5 6485.001125625626u,0 6488.910285785786u,0 6488.911285785786u,1.5 6490.865365865866u,1.5 6490.866365865866u,0 6496.730606106106u,0 6496.7316061061065u,1.5 6497.708146146146u,1.5 6497.709146146146u,0 6500.640766266267u,0 6500.641766266267u,1.5 6501.618306306306u,1.5 6501.6193063063065u,0 6511.393706706706u,0 6511.3947067067065u,1.5 6512.371246746747u,1.5 6512.372246746747u,0 6513.348786786787u,0 6513.349786786787u,1.5 6514.3263268268265u,1.5 6514.327326826827u,0 6517.258946946947u,0 6517.259946946947u,1.5 6518.236486986987u,1.5 6518.237486986987u,0 6520.191567067067u,0 6520.192567067067u,1.5 6521.169107107107u,1.5 6521.1701071071075u,0 6525.079267267268u,0 6525.080267267268u,1.5 6527.034347347347u,1.5 6527.035347347347u,0 6528.9894274274275u,0 6528.990427427428u,1.5 6532.899587587588u,1.5 6532.900587587588u,0 6533.8771276276275u,0 6533.878127627628u,1.5 6535.832207707707u,1.5 6535.8332077077075u,0 6536.809747747748u,0 6536.810747747748u,1.5 6543.6525280280275u,1.5 6543.653528028028u,0 6544.630068068068u,0 6544.631068068068u,1.5 6549.517768268269u,1.5 6549.518768268269u,0 6551.472848348348u,0 6551.473848348348u,1.5 6553.4279284284285u,1.5 6553.428928428429u,0 6562.225788788789u,0 6562.226788788789u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6565.158408908908u,1.5 6565.1594089089085u,0 6566.135948948949u,0 6566.136948948949u,1.5 6568.0910290290285u,1.5 6568.092029029029u,0 6569.068569069069u,0 6569.069569069069u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.001189189189u,0 6572.002189189189u,1.5 6574.933809309309u,1.5 6574.9348093093095u,0 6575.911349349349u,0 6575.912349349349u,1.5 6577.866429429429u,1.5 6577.86742942943u,0 6586.66428978979u,0 6586.66528978979u,1.5 6587.6418298298295u,1.5 6587.64282982983u,0 6588.61936986987u,0 6588.62036986987u,1.5 6590.57444994995u,1.5 6590.57544994995u,0 6592.5295300300295u,0 6592.53053003003u,1.5 6596.43969019019u,1.5 6596.44069019019u,0 6597.4172302302295u,0 6597.41823023023u,1.5 6598.394770270271u,1.5 6598.395770270271u,0 6600.34985035035u,0 6600.35085035035u,1.5 6601.32739039039u,1.5 6601.32839039039u,0 6602.30493043043u,0 6602.305930430431u,1.5 6603.282470470471u,1.5 6603.283470470471u,0 6604.26001051051u,0 6604.2610105105105u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6607.19263063063u,0 6607.193630630631u,1.5 6612.0803308308305u,1.5 6612.081330830831u,0 6613.057870870871u,0 6613.058870870871u,1.5 6614.03541091091u,1.5 6614.0364109109105u,0 6615.012950950951u,0 6615.013950950951u,1.5 6615.990490990991u,1.5 6615.991490990991u,0 6617.945571071071u,0 6617.946571071071u,1.5 6619.900651151151u,1.5 6619.901651151151u,0 6621.8557312312305u,0 6621.856731231231u,1.5 6623.810811311311u,1.5 6623.811811311311u,0 6624.788351351351u,0 6624.789351351351u,1.5 6626.743431431431u,1.5 6626.744431431432u,0 6627.720971471472u,0 6627.721971471472u,1.5 6629.676051551551u,1.5 6629.677051551551u,0 6631.631131631631u,0 6631.632131631632u,1.5 6632.608671671672u,1.5 6632.609671671672u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6637.496371871872u,0 6637.497371871872u,1.5 6638.473911911911u,1.5 6638.4749119119115u,0 6639.451451951952u,0 6639.452451951952u,1.5 6643.361612112112u,1.5 6643.362612112112u,0 6645.316692192192u,0 6645.317692192192u,1.5 6646.2942322322315u,1.5 6646.295232232232u,0 6649.226852352352u,0 6649.227852352352u,1.5 6650.204392392392u,1.5 6650.205392392392u,0 6651.181932432432u,0 6651.182932432433u,1.5 6654.114552552552u,1.5 6654.115552552552u,0 6655.092092592593u,0 6655.093092592593u,1.5 6657.047172672673u,1.5 6657.048172672673u,0 6659.002252752753u,0 6659.003252752753u,1.5 6659.979792792793u,1.5 6659.980792792793u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6664.867492992993u,1.5 6664.868492992993u,0 6666.822573073073u,0 6666.823573073073u,1.5 6668.777653153153u,1.5 6668.778653153153u,0 6672.687813313313u,0 6672.688813313313u,1.5 6673.665353353353u,1.5 6673.666353353353u,0 6674.642893393393u,0 6674.643893393393u,1.5 6676.597973473474u,1.5 6676.598973473474u,0 6677.575513513513u,0 6677.576513513513u,1.5 6678.553053553553u,1.5 6678.554053553553u,0 6679.530593593594u,0 6679.531593593594u,1.5 6680.508133633633u,1.5 6680.509133633634u,0 6684.418293793794u,0 6684.419293793794u,1.5 6691.261074074074u,1.5 6691.262074074074u,0 6693.216154154154u,0 6693.217154154154u,1.5 6694.193694194194u,1.5 6694.194694194194u,0 6698.103854354354u,0 6698.104854354354u,1.5 6702.991554554554u,1.5 6702.992554554554u,0 6704.946634634634u,0 6704.947634634635u,1.5 6706.901714714714u,1.5 6706.902714714714u,0 6707.879254754755u,0 6707.880254754755u,1.5 6708.856794794795u,1.5 6708.857794794795u,0 6709.834334834834u,0 6709.835334834835u,1.5 6711.789414914914u,1.5 6711.790414914914u,0 6712.766954954955u,0 6712.767954954955u,1.5 6713.744494994995u,1.5 6713.745494994995u,0 6715.699575075075u,0 6715.700575075075u,1.5 6716.677115115115u,1.5 6716.678115115115u,0 6718.632195195195u,0 6718.633195195195u,1.5 6719.609735235234u,1.5 6719.610735235235u,0 6720.587275275276u,0 6720.588275275276u,1.5 6723.519895395395u,1.5 6723.520895395395u,0 6726.452515515515u,0 6726.453515515515u,1.5 6727.430055555555u,1.5 6727.431055555555u,0 6729.385135635635u,0 6729.386135635636u,1.5 6733.295295795796u,1.5 6733.296295795796u,0 6734.272835835835u,0 6734.273835835836u,1.5 6735.250375875876u,1.5 6735.251375875876u,0 6736.227915915916u,0 6736.228915915916u,1.5 6737.205455955956u,1.5 6737.206455955956u,0 6741.115616116116u,0 6741.116616116116u,1.5 6742.093156156156u,1.5 6742.094156156156u,0 6743.070696196196u,0 6743.071696196196u,1.5 6744.048236236235u,1.5 6744.049236236236u,0 6745.025776276277u,0 6745.026776276277u,1.5 6746.003316316316u,1.5 6746.004316316316u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6753.823636636636u,0 6753.824636636637u,1.5 6754.801176676677u,1.5 6754.802176676677u,0 6761.6439569569575u,0 6761.644956956958u,1.5 6766.5316571571575u,1.5 6766.532657157158u,0 6768.486737237236u,0 6768.487737237237u,1.5 6769.464277277278u,1.5 6769.465277277278u,0 6771.4193573573575u,0 6771.420357357358u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6775.329517517517u,1.5 6775.330517517517u,0 6776.3070575575575u,0 6776.308057557558u,1.5 6777.284597597598u,1.5 6777.285597597598u,0 6778.262137637637u,0 6778.263137637638u,1.5 6779.239677677678u,1.5 6779.240677677678u,0 6780.217217717717u,0 6780.218217717717u,1.5 6782.172297797798u,1.5 6782.173297797798u,0 6783.149837837837u,0 6783.150837837838u,1.5 6786.0824579579585u,1.5 6786.083457957959u,0 6787.059997997998u,0 6787.060997997998u,1.5 6788.037538038037u,1.5 6788.038538038038u,0 6791.947698198198u,0 6791.948698198198u,1.5 6794.880318318318u,1.5 6794.881318318318u,0 6795.8578583583585u,0 6795.858858358359u,1.5 6798.790478478479u,1.5 6798.791478478479u,0 6802.700638638638u,0 6802.7016386386385u,1.5 6803.678178678679u,1.5 6803.679178678679u,0 6805.633258758759u,0 6805.63425875876u,1.5 6808.565878878879u,1.5 6808.566878878879u,0 6810.520958958959u,0 6810.52195895896u,1.5 6811.498498998999u,1.5 6811.499498998999u,0 6813.453579079079u,0 6813.454579079079u,1.5 6814.431119119119u,1.5 6814.432119119119u,0 6815.4086591591595u,0 6815.40965915916u,1.5 6818.34127927928u,1.5 6818.34227927928u,0 6819.318819319319u,0 6819.319819319319u,1.5 6821.273899399399u,1.5 6821.274899399399u,0 6823.22897947948u,0 6823.22997947948u,1.5 6824.206519519519u,1.5 6824.207519519519u,0 6826.1615995996u,0 6826.1625995996u,1.5 6827.139139639639u,1.5 6827.1401396396395u,0 6828.11667967968u,0 6828.11767967968u,1.5 6831.0492997998u,1.5 6831.0502997998u,0 6832.026839839839u,0 6832.0278398398395u,1.5 6833.00437987988u,1.5 6833.00537987988u,0 6833.98191991992u,0 6833.98291991992u,1.5 6834.95945995996u,1.5 6834.960459959961u,0 6835.937u,0 6835.938u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6839.8471601601605u,0 6839.848160160161u,1.5 6841.802240240239u,1.5 6841.80324024024u,0 6842.779780280281u,0 6842.780780280281u,1.5 6844.7348603603605u,1.5 6844.735860360361u,0 6845.7124004004u,0 6845.7134004004u,1.5 6846.68994044044u,1.5 6846.6909404404405u,0 6848.64502052052u,0 6848.64602052052u,1.5 6849.6225605605605u,1.5 6849.623560560561u,0 6851.57764064064u,0 6851.5786406406405u,1.5 6854.510260760761u,1.5 6854.511260760762u,0 6856.46534084084u,0 6856.4663408408405u,1.5 6857.442880880881u,1.5 6857.443880880881u,0 6859.397960960961u,0 6859.398960960962u,1.5 6861.35304104104u,1.5 6861.354041041041u,0 6864.285661161161u,0 6864.286661161162u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6867.218281281282u,0 6867.219281281282u,1.5 6870.150901401401u,1.5 6870.151901401401u,0 6871.128441441441u,0 6871.1294414414415u,1.5 6872.105981481482u,1.5 6872.106981481482u,0 6876.016141641641u,0 6876.0171416416415u,1.5 6876.993681681682u,1.5 6876.994681681682u,0 6878.948761761762u,0 6878.949761761763u,1.5 6884.814002002002u,1.5 6884.815002002002u,0 6885.791542042041u,0 6885.7925420420415u,1.5 6886.769082082082u,1.5 6886.770082082082u,0 6892.634322322322u,0 6892.635322322322u,1.5 6893.611862362362u,1.5 6893.612862362363u,0 6896.544482482483u,0 6896.545482482483u,1.5 6900.454642642642u,1.5 6900.4556426426425u,0 6901.432182682683u,0 6901.433182682683u,1.5 6903.387262762763u,1.5 6903.388262762764u,0 6907.297422922923u,0 6907.298422922923u,1.5 6909.252503003003u,1.5 6909.253503003003u,0 6912.185123123123u,0 6912.186123123123u,1.5 6913.162663163163u,1.5 6913.163663163164u,0 6914.140203203203u,0 6914.141203203203u,1.5 6920.982983483484u,1.5 6920.983983483484u,0 6922.938063563563u,0 6922.939063563564u,1.5 6924.893143643643u,1.5 6924.8941436436435u,0 6926.848223723723u,0 6926.849223723723u,1.5 6927.825763763764u,1.5 6927.826763763765u,0 6932.713463963964u,0 6932.714463963965u,1.5 6933.691004004004u,1.5 6933.692004004004u,0 6934.668544044043u,0 6934.6695440440435u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6936.623624124124u,0 6936.624624124124u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6939.556244244243u,0 6939.5572442442435u,1.5 6942.488864364364u,1.5 6942.489864364365u,0 6943.466404404404u,0 6943.467404404404u,1.5 6945.421484484485u,1.5 6945.422484484485u,0 6946.399024524524u,0 6946.400024524524u,1.5 6950.309184684685u,1.5 6950.310184684685u,0 6954.219344844844u,0 6954.2203448448445u,1.5 6955.196884884885u,1.5 6955.197884884885u,0 6958.129505005005u,0 6958.130505005005u,1.5 6959.107045045044u,1.5 6959.1080450450445u,0 6962.039665165165u,0 6962.040665165166u,1.5 6963.017205205205u,1.5 6963.018205205205u,0 6963.994745245244u,0 6963.9957452452445u,1.5 6964.972285285286u,1.5 6964.973285285286u,0 6967.904905405405u,0 6967.905905405405u,1.5 6968.882445445445u,1.5 6968.883445445445u,0 6969.859985485486u,0 6969.860985485486u,1.5 6970.837525525525u,1.5 6970.838525525525u,0 6971.815065565565u,0 6971.816065565566u,1.5 6972.792605605606u,1.5 6972.793605605606u,0 6973.770145645645u,0 6973.771145645645u,1.5 6974.747685685686u,1.5 6974.748685685686u,0 6976.702765765766u,0 6976.703765765767u,1.5 6978.657845845845u,1.5 6978.6588458458455u,0 6980.612925925926u,0 6980.613925925926u,1.5 6981.590465965966u,1.5 6981.591465965967u,0 6982.568006006006u,0 6982.569006006006u,1.5 6986.478166166166u,1.5 6986.479166166167u,0 6987.455706206206u,0 6987.456706206206u,1.5 6988.433246246245u,1.5 6988.4342462462455u,0 6990.388326326326u,0 6990.389326326326u,1.5 6991.365866366366u,1.5 6991.366866366367u,0 6992.343406406406u,0 6992.344406406406u,1.5 6994.298486486487u,1.5 6994.299486486487u,0 6995.276026526526u,0 6995.277026526526u,1.5
vb12 b12 0 pwl 0,0  3.90966016016016u,0 3.9106601601601603u,1.5 4.8872002002002u,1.5 4.8882002002002u,0 10.75244044044044u,0 10.753440440440441u,1.5 11.72998048048048u,1.5 11.730980480480481u,0 12.70752052052052u,0 12.708520520520521u,1.5 13.68506056056056u,1.5 13.686060560560561u,0 17.59522072072072u,0 17.59622072072072u,1.5 18.572760760760765u,1.5 18.573760760760763u,0 25.415541041041042u,0 25.41654104104104u,1.5 26.393081081081085u,1.5 26.394081081081083u,0 27.370621121121122u,0 27.37162112112112u,1.5 28.348161161161162u,1.5 28.34916116116116u,0 30.303241241241246u,0 30.304241241241243u,1.5 31.280781281281282u,1.5 31.28178128128128u,0 33.23586136136136u,0 33.23686136136136u,1.5 35.19094144144144u,1.5 35.19194144144144u,0 36.16848148148148u,0 36.16948148148148u,1.5 37.146021521521526u,1.5 37.14702152152153u,0 38.12356156156156u,0 38.12456156156156u,1.5 40.07864164164164u,1.5 40.07964164164164u,0 41.05618168168168u,0 41.05718168168168u,1.5 58.6519024024024u,1.5 58.652902402402404u,0 59.62944244244244u,0 59.630442442442444u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 85.04548348348348u,0 85.04648348348348u,1.5 86.02302352352352u,1.5 86.02402352352352u,0 87.00056356356356u,0 87.00156356356356u,1.5 90.91072372372372u,1.5 90.91172372372372u,0 91.88826376376376u,0 91.88926376376376u,1.5 104.59628428428428u,1.5 104.59728428428429u,0 106.55136436436436u,0 106.55236436436437u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 109.48398448448448u,0 109.48498448448449u,1.5 110.46152452452452u,1.5 110.46252452452453u,0 116.32676476476476u,0 116.32776476476477u,1.5 117.3043048048048u,1.5 117.3053048048048u,0 123.16954504504503u,0 123.17054504504503u,1.5 124.14708508508508u,1.5 124.14808508508509u,0 125.12462512512512u,0 125.12562512512513u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 136.85510560560562u,0 136.8561056056056u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 150.54066616616618u,0 150.54166616616615u,1.5 152.49574624624626u,1.5 152.49674624624623u,0 153.4732862862863u,0 153.4742862862863u,1.5 158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 164.22622672672674u,1.5 164.2272267267267u,0 174.97916716716716u,0 174.98016716716714u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 185.73210760760762u,0 185.7331076076076u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 188.66472772772775u,1.5 188.66572772772773u,0 195.50750800800802u,0 195.508508008008u,1.5 197.4625880880881u,1.5 197.46358808808807u,0 198.44012812812815u,0 198.44112812812813u,1.5 207.2379884884885u,1.5 207.23898848848847u,0 208.21552852852852u,0 208.2165285285285u,1.5 210.17060860860863u,1.5 210.1716086086086u,0 218.96846896896898u,0 218.96946896896895u,1.5 219.94600900900903u,1.5 219.947009009009u,0 220.92354904904906u,0 220.92454904904903u,1.5 229.72140940940943u,1.5 229.7224094094094u,0 230.69894944944946u,0 230.69994944944943u,1.5 231.6764894894895u,1.5 231.6774894894895u,0 237.54172972972972u,0 237.5427297297297u,1.5 238.51926976976978u,1.5 238.52026976976975u,0 239.4968098098098u,0 239.49780980980978u,1.5 240.47434984984986u,1.5 240.47534984984983u,0 241.4518898898899u,0 241.4528898898899u,1.5 242.42942992992997u,1.5 242.43042992992994u,0 243.40696996996996u,0 243.40796996996994u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 259.04761061061066u,0 259.04861061061064u,1.5 260.02515065065063u,1.5 260.0261506506506u,0 261.00269069069066u,0 261.00369069069063u,1.5 261.98023073073074u,1.5 261.9812307307307u,0 262.95777077077076u,0 262.95877077077074u,1.5 270.77809109109114u,1.5 270.7790910910911u,0 271.75563113113117u,0 271.75663113113114u,1.5 272.73317117117114u,1.5 272.7341711711711u,0 279.57595145145143u,0 279.5769514514514u,1.5 280.5534914914915u,1.5 280.5544914914915u,0 281.53103153153154u,0 281.5320315315315u,1.5 282.50857157157157u,1.5 282.50957157157154u,0 283.48611161161165u,0 283.4871116116116u,1.5 289.35135185185186u,1.5 289.35235185185184u,0 290.32889189189194u,0 290.3298918918919u,1.5 294.23905205205205u,1.5 294.240052052052u,0 302.0593723723724u,0 302.0603723723724u,1.5 304.0144524524524u,1.5 304.0154524524524u,0 305.9695325325325u,0 305.9705325325325u,1.5 306.9470725725726u,1.5 306.9480725725726u,0 307.92461261261263u,0 307.9256126126126u,1.5 313.78985285285285u,1.5 313.7908528528528u,0 314.76739289289293u,0 314.7683928928929u,1.5 315.74493293293295u,1.5 315.74593293293293u,0 317.700013013013u,0 317.701013013013u,1.5 318.67755305305303u,1.5 318.678553053053u,0 323.5652532532532u,0 323.5662532532532u,1.5 324.5427932932933u,1.5 324.5437932932933u,0 326.4978733733734u,0 326.4988733733734u,1.5 328.45295345345346u,1.5 328.45395345345344u,0 329.4304934934935u,0 329.43149349349346u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 336.2732737737738u,0 336.27427377377376u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 338.2283538538539u,0 338.22935385385387u,1.5 340.18343393393394u,1.5 340.1844339339339u,0 349.9588343343343u,0 349.9598343343343u,1.5 350.9363743743744u,1.5 350.9373743743744u,0 351.9139144144144u,0 351.9149144144144u,1.5 352.8914544544545u,1.5 352.8924544544545u,0 353.8689944944945u,0 353.86999449449445u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 374.39733533533536u,0 374.39833533533533u,1.5 375.3748753753754u,1.5 375.37587537537536u,0 378.3074954954955u,0 378.3084954954955u,1.5 380.26257557557557u,1.5 380.26357557557554u,0 381.2401156156156u,0 381.24111561561557u,1.5 389.06043593593597u,1.5 389.06143593593595u,0 390.037975975976u,0 390.038975975976u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 395.90321621621626u,1.5 395.90421621621624u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 405.67861661661664u,0 405.6796166166166u,1.5 406.65615665665666u,1.5 406.65715665665664u,0 408.61123673673677u,0 408.61223673673675u,1.5 409.5887767767768u,1.5 409.5897767767768u,0 410.5663168168168u,0 410.5673168168168u,1.5 411.54385685685685u,1.5 411.5448568568568u,0 412.5213968968969u,0 412.52239689689685u,1.5 414.476476976977u,1.5 414.47747697697696u,0 415.45401701701707u,0 415.45501701701704u,1.5 432.07219769769773u,1.5 432.0731976976977u,0 433.04973773773776u,0 433.05073773773773u,1.5 434.0272777777778u,1.5 434.02827777777776u,0 435.00481781781787u,0 435.00581781781784u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 437.93743793793794u,0 437.9384379379379u,1.5 438.91497797797797u,1.5 438.91597797797795u,0 455.53315865865864u,0 455.5341586586586u,1.5 456.5106986986987u,1.5 456.5116986986987u,0 462.37593893893893u,0 462.3769389389389u,1.5 463.353478978979u,1.5 463.354478978979u,0 466.28609909909915u,0 466.2870990990991u,1.5 468.2411791791792u,1.5 468.2421791791792u,0 470.19625925925925u,0 470.1972592592592u,1.5 471.17379929929933u,1.5 471.1747992992993u,0 472.15133933933936u,0 472.15233933933933u,1.5 474.1064194194194u,1.5 474.1074194194194u,0 475.08395945945944u,0 475.0849594594594u,1.5 476.0614994994995u,1.5 476.0624994994995u,0 478.0165795795796u,0 478.0175795795796u,1.5 486.8144399399399u,1.5 486.8154399399399u,0 487.79197997998u,0 487.79297997998u,1.5 488.7695200200201u,1.5 488.77052002002006u,0 489.7470600600601u,0 489.7480600600601u,1.5 496.58984034034034u,1.5 496.5908403403403u,0 497.56738038038037u,0 497.56838038038035u,1.5 503.4326206206207u,1.5 503.4336206206207u,0 504.41016066066067u,0 504.41116066066064u,1.5 509.2978608608609u,1.5 509.2988608608609u,0 510.2754009009009u,0 510.27640090090085u,1.5 518.0957212212213u,1.5 518.0967212212213u,0 519.0732612612613u,0 519.0742612612613u,1.5 521.0283413413413u,1.5 521.0293413413413u,0 522.0058813813813u,0 522.0068813813813u,1.5 525.9160415415415u,1.5 525.9170415415415u,0 526.8935815815815u,0 526.8945815815815u,1.5 528.8486616616617u,1.5 528.8496616616617u,0 530.8037417417418u,0 530.8047417417417u,1.5 531.7812817817818u,1.5 531.7822817817818u,0 533.7363618618618u,0 533.7373618618618u,1.5 534.7139019019019u,1.5 534.7149019019018u,0 540.5791421421421u,0 540.5801421421421u,1.5 541.5566821821823u,1.5 541.5576821821822u,0 560.1299429429429u,0 560.1309429429429u,1.5 561.107482982983u,1.5 561.108482982983u,0 563.0625630630631u,0 563.063563063063u,1.5 564.0401031031031u,1.5 564.0411031031031u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 569.9053433433434u,0 569.9063433433433u,1.5 584.5684439439439u,1.5 584.5694439439438u,0 585.545983983984u,0 585.546983983984u,1.5 587.501064064064u,1.5 587.502064064064u,0 589.4561441441441u,0 589.4571441441441u,1.5 590.4336841841842u,1.5 590.4346841841842u,0 592.3887642642643u,0 592.3897642642643u,1.5 593.3663043043043u,1.5 593.3673043043043u,0 596.2989244244244u,0 596.2999244244244u,1.5 597.2764644644644u,1.5 597.2774644644644u,0 602.1641646646647u,0 602.1651646646646u,1.5 603.1417047047047u,1.5 603.1427047047047u,0 605.0967847847849u,0 605.0977847847848u,1.5 606.0743248248249u,1.5 606.0753248248249u,0 607.0518648648649u,0 607.0528648648649u,1.5 620.7374254254254u,1.5 620.7384254254254u,0 621.7149654654654u,0 621.7159654654654u,1.5 623.6700455455456u,1.5 623.6710455455456u,0 637.355606106106u,0 637.356606106106u,1.5 649.0860865865866u,1.5 649.0870865865866u,0 660.816567067067u,0 660.817567067067u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 662.7716471471472u,0 662.7726471471472u,1.5 663.7491871871872u,1.5 663.7501871871872u,0 664.7267272272272u,0 664.7277272272272u,1.5 672.5470475475475u,1.5 672.5480475475475u,0 674.5021276276276u,0 674.5031276276276u,1.5 675.4796676676676u,1.5 675.4806676676676u,0 685.255068068068u,0 685.256068068068u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 696.0080085085085u,1.5 696.0090085085085u,0 696.9855485485485u,0 696.9865485485485u,1.5 697.9630885885886u,1.5 697.9640885885885u,0 707.7384889889889u,0 707.7394889889889u,1.5 708.716029029029u,1.5 708.7170290290289u,0 709.693569069069u,0 709.694569069069u,1.5 716.5363493493494u,1.5 716.5373493493494u,0 717.5138893893894u,0 717.5148893893894u,1.5 718.4914294294294u,1.5 718.4924294294294u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 729.24436986987u,0 729.2453698698699u,1.5 730.22190990991u,1.5 730.22290990991u,0 731.19944994995u,0 731.20044994995u,1.5 739.0197702702703u,1.5 739.0207702702703u,0 740.9748503503504u,0 740.9758503503504u,1.5 741.9523903903904u,1.5 741.9533903903904u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 761.5031911911911u,1.5 761.5041911911911u,0 762.4807312312312u,0 762.4817312312312u,1.5 763.4582712712713u,1.5 763.4592712712713u,0 770.3010515515515u,0 770.3020515515515u,1.5 771.2785915915915u,1.5 771.2795915915915u,0 772.2561316316315u,0 772.2571316316315u,1.5 781.053991991992u,1.5 781.054991991992u,0 782.031532032032u,0 782.032532032032u,1.5 783.0090720720721u,1.5 783.010072072072u,0 790.8293923923924u,0 790.8303923923924u,1.5 792.7844724724725u,1.5 792.7854724724725u,0 793.7620125125126u,0 793.7630125125125u,1.5 803.5374129129129u,1.5 803.5384129129129u,0 814.2903533533533u,0 814.2913533533533u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 816.2454334334335u,0 816.2464334334335u,1.5 825.0432937937937u,1.5 825.0442937937937u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 841.6614744744745u,0 841.6624744744745u,1.5 848.5042547547547u,1.5 848.5052547547547u,0 849.4817947947948u,0 849.4827947947948u,1.5 851.4368748748749u,1.5 851.4378748748749u,0 854.3694949949951u,0 854.370494994995u,1.5 855.3470350350351u,1.5 855.3480350350351u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 868.0550555555556u,1.5 868.0560555555555u,0 869.0325955955957u,0 869.0335955955957u,1.5 878.8079959959961u,1.5 878.808995995996u,0 894.4486366366367u,0 894.4496366366367u,1.5 896.4037167167166u,1.5 896.4047167167166u,0 897.3812567567567u,0 897.3822567567566u,1.5 908.1341971971972u,1.5 908.1351971971972u,0 909.1117372372372u,0 909.1127372372372u,1.5 911.0668173173173u,1.5 911.0678173173172u,0 912.0443573573574u,0 912.0453573573574u,1.5 913.0218973973974u,1.5 913.0228973973974u,0 913.9994374374375u,0 914.0004374374374u,1.5 914.9769774774775u,1.5 914.9779774774775u,0 916.9320575575576u,0 916.9330575575576u,1.5 917.9095975975977u,1.5 917.9105975975976u,0 927.684997997998u,0 927.685997997998u,1.5 928.6625380380381u,1.5 928.663538038038u,0 932.5726981981983u,0 932.5736981981983u,1.5 933.5502382382382u,1.5 933.5512382382382u,0 935.5053183183182u,0 935.5063183183182u,1.5 938.4379384384384u,1.5 938.4389384384384u,0 939.4154784784785u,0 939.4164784784784u,1.5 959.9438193193192u,1.5 959.9448193193192u,0 960.9213593593594u,0 960.9223593593593u,1.5 964.8315195195195u,1.5 964.8325195195195u,0 966.7865995995996u,0 966.7875995995996u,1.5 967.7641396396397u,1.5 967.7651396396396u,0 968.7416796796797u,0 968.7426796796797u,1.5 970.6967597597597u,1.5 970.6977597597597u,0 972.6518398398398u,0 972.6528398398398u,1.5 973.6293798798798u,1.5 973.6303798798798u,0 974.60691991992u,0 974.6079199199199u,1.5 975.58445995996u,1.5 975.58545995996u,0 977.5395400400402u,0 977.5405400400401u,1.5 978.5170800800801u,1.5 978.51808008008u,0 981.4497002002003u,0 981.4507002002002u,1.5 982.4272402402403u,1.5 982.4282402402403u,0 983.4047802802802u,0 983.4057802802802u,1.5 984.3823203203203u,1.5 984.3833203203203u,0 989.2700205205206u,0 989.2710205205206u,1.5 990.2475605605605u,1.5 990.2485605605605u,0 991.2251006006006u,0 991.2261006006006u,1.5 992.2026406406408u,1.5 992.2036406406407u,0 994.1577207207208u,0 994.1587207207208u,1.5 995.1352607607607u,1.5 995.1362607607607u,0 999.045420920921u,0 999.0464209209209u,1.5 1000.0229609609609u,1.5 1000.0239609609608u,0 1001.9780410410411u,0 1001.9790410410411u,1.5 1002.955581081081u,1.5 1002.956581081081u,0 1004.9106611611611u,0 1004.9116611611611u,1.5 1005.8882012012012u,1.5 1005.8892012012012u,0 1013.7085215215216u,0 1013.7095215215215u,1.5 1014.6860615615615u,1.5 1014.6870615615614u,0 1016.6411416416418u,0 1016.6421416416417u,1.5 1017.6186816816817u,1.5 1017.6196816816816u,0 1021.5288418418419u,0 1021.5298418418419u,1.5 1022.5063818818818u,1.5 1022.5073818818818u,0 1026.416542042042u,0 1026.4175420420422u,1.5 1027.394082082082u,1.5 1027.3950820820821u,0 1028.371622122122u,0 1028.3726221221223u,1.5 1029.349162162162u,1.5 1029.3501621621622u,0 1030.3267022022021u,0 1030.3277022022023u,1.5 1031.3042422422423u,1.5 1031.3052422422425u,0 1032.2817822822822u,0 1032.2827822822824u,1.5 1033.2593223223223u,1.5 1033.2603223223225u,0 1034.2368623623622u,0 1034.2378623623624u,1.5 1057.6978233233233u,1.5 1057.6988233233235u,0 1058.6753633633632u,0 1058.6763633633634u,1.5 1061.6079834834834u,1.5 1061.6089834834836u,0 1062.5855235235235u,0 1062.5865235235237u,1.5 1065.5181436436435u,1.5 1065.5191436436437u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1070.4058438438437u,0 1070.406843843844u,1.5 1071.3833838838837u,1.5 1071.3843838838839u,0 1086.0464844844844u,0 1086.0474844844846u,1.5 1087.0240245245245u,1.5 1087.0250245245247u,0 1088.9791046046046u,0 1088.9801046046048u,1.5 1089.9566446446445u,1.5 1089.9576446446447u,0 1091.9117247247245u,0 1091.9127247247247u,1.5 1092.8892647647647u,1.5 1092.8902647647649u,0 1093.8668048048046u,0 1093.8678048048048u,1.5 1102.6646651651652u,1.5 1102.6656651651654u,0 1103.642205205205u,0 1103.6432052052053u,1.5 1104.6197452452452u,1.5 1104.6207452452454u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1107.5523653653654u,1.5 1107.5533653653656u,0 1108.5299054054053u,0 1108.5309054054055u,1.5 1109.5074454454455u,1.5 1109.5084454454457u,0 1120.2603858858856u,0 1120.2613858858858u,1.5 1121.2379259259258u,1.5 1121.238925925926u,0 1122.215465965966u,0 1122.216465965966u,1.5 1124.170546046046u,1.5 1124.1715460460462u,0 1125.1480860860859u,0 1125.149086086086u,1.5 1134.9234864864864u,1.5 1134.9244864864866u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1148.609047047047u,0 1148.6100470470471u,1.5 1150.564127127127u,1.5 1150.5651271271272u,0 1151.5416671671671u,0 1151.5426671671673u,1.5 1152.519207207207u,1.5 1152.5202072072072u,0 1153.4967472472472u,0 1153.4977472472474u,1.5 1154.474287287287u,1.5 1154.4752872872873u,0 1155.4518273273272u,0 1155.4528273273274u,1.5 1161.3170675675676u,1.5 1161.3180675675678u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1163.2721476476477u,1.5 1163.2731476476479u,0 1164.2496876876876u,0 1164.2506876876878u,1.5 1165.2272277277275u,1.5 1165.2282277277277u,0 1172.0700080080078u,0 1172.071008008008u,1.5 1173.047548048048u,1.5 1173.0485480480481u,0 1175.002628128128u,0 1175.0036281281282u,1.5 1177.9352482482482u,1.5 1177.9362482482484u,0 1178.912788288288u,0 1178.9137882882883u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1197.486049049049u,0 1197.4870490490491u,1.5 1199.441129129129u,1.5 1199.4421291291292u,0 1200.418669169169u,0 1200.4196691691693u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1208.2389894894895u,0 1208.2399894894897u,1.5 1210.1940695695696u,1.5 1210.1950695695698u,0 1217.0368498498497u,0 1217.0378498498499u,1.5 1218.0143898898898u,1.5 1218.01538988989u,0 1218.9919299299297u,0 1218.99292992993u,1.5 1219.9694699699699u,1.5 1219.97046996997u,0 1220.9470100100098u,0 1220.94801001001u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1231.6999504504504u,1.5 1231.7009504504506u,0 1241.4753508508506u,0 1241.4763508508508u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1254.1833713713713u,1.5 1254.1843713713715u,0 1260.0486116116115u,0 1260.0496116116117u,1.5 1261.0261516516516u,1.5 1261.0271516516518u,0 1262.0036916916918u,0 1262.004691691692u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1269.8240120120117u,0 1269.825012012012u,1.5 1270.8015520520519u,1.5 1270.802552052052u,0 1271.779092092092u,0 1271.7800920920922u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1280.5769524524524u,0 1280.5779524524526u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1291.3298928928928u,0 1291.330892892893u,1.5 1292.3074329329327u,1.5 1292.3084329329329u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1303.0603733733733u,0 1303.0613733733735u,1.5 1305.0154534534533u,1.5 1305.0164534534536u,0 1305.9929934934935u,0 1305.9939934934937u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1315.7683938938937u,0 1315.769393893894u,1.5 1316.7459339339337u,1.5 1316.7469339339339u,0 1327.4988743743743u,0 1327.4998743743745u,1.5 1329.4539544544543u,1.5 1329.4549544544545u,0 1330.4314944944945u,0 1330.4324944944947u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1342.1619749749748u,1.5 1342.162974974975u,0 1348.0272152152152u,0 1348.0282152152154u,1.5 1349.004755255255u,1.5 1349.0057552552553u,0 1350.9598353353351u,0 1350.9608353353353u,1.5 1352.9149154154154u,1.5 1352.9159154154156u,0 1353.8924554554553u,0 1353.8934554554555u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1367.578016016016u,0 1367.579016016016u,1.5 1368.5555560560558u,1.5 1368.556556056056u,0 1376.3758763763763u,0 1376.3768763763765u,1.5 1377.3534164164164u,1.5 1377.3544164164166u,0 1378.3309564564563u,0 1378.3319564564565u,1.5 1379.3084964964964u,1.5 1379.3094964964966u,0 1380.2860365365364u,0 1380.2870365365366u,1.5 1384.1961966966967u,1.5 1384.197196696697u,0 1385.1737367367366u,0 1385.1747367367368u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1400.8143773773772u,0 1400.8153773773774u,1.5 1401.7919174174174u,1.5 1401.7929174174176u,0 1408.6346976976977u,0 1408.6356976976979u,1.5 1409.6122377377376u,1.5 1409.6132377377378u,0 1411.5673178178179u,0 1411.568317817818u,1.5 1414.4999379379378u,1.5 1414.500937937938u,0 1415.4774779779777u,0 1415.478477977978u,1.5 1431.1181186186186u,1.5 1431.1191186186188u,0 1432.0956586586585u,0 1432.0966586586587u,1.5 1433.0731986986987u,1.5 1433.0741986986989u,0 1434.0507387387386u,0 1434.0517387387388u,1.5 1436.0058188188189u,1.5 1436.006818818819u,0 1438.938438938939u,0 1438.9394389389392u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1464.35447997998u,0 1464.3554799799801u,1.5 1465.3320200200199u,1.5 1465.33302002002u,0 1467.2871001001u,0 1467.2881001001u,1.5 1468.26464014014u,1.5 1468.2656401401402u,0 1470.21972022022u,0 1470.2207202202203u,1.5 1471.19726026026u,1.5 1471.1982602602602u,0 1473.1523403403403u,0 1473.1533403403405u,1.5 1474.1298803803802u,1.5 1474.1308803803804u,0 1476.0849604604603u,0 1476.0859604604605u,1.5 1477.0625005005004u,1.5 1477.0635005005006u,0 1478.0400405405405u,0 1478.0410405405407u,1.5 1480.9726606606605u,1.5 1480.9736606606607u,0 1481.9502007007006u,0 1481.9512007007008u,1.5 1482.9277407407408u,1.5 1482.928740740741u,0 1483.9052807807807u,0 1483.906280780781u,1.5 1494.658221221221u,1.5 1494.6592212212213u,0 1495.635761261261u,0 1495.6367612612612u,1.5 1513.231481981982u,1.5 1513.2324819819821u,0 1514.209022022022u,0 1514.2100220220223u,1.5 1520.074262262262u,1.5 1520.0752622622622u,0 1521.0518023023021u,0 1521.0528023023023u,1.5 1522.0293423423423u,1.5 1522.0303423423425u,0 1523.0068823823822u,0 1523.0078823823824u,1.5 1524.9619624624622u,1.5 1524.9629624624624u,0 1525.9395025025024u,0 1525.9405025025026u,1.5 1526.9170425425425u,1.5 1526.9180425425427u,0 1527.8945825825824u,0 1527.8955825825826u,1.5 1530.8272027027026u,1.5 1530.8282027027028u,0 1531.8047427427427u,0 1531.805742742743u,1.5 1532.7822827827827u,1.5 1532.7832827827829u,0 1562.108483983984u,0 1562.109483983984u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1565.041104104104u,0 1565.0421041041043u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1567.973724224224u,0 1567.9747242242242u,1.5 1579.7042047047046u,1.5 1579.7052047047048u,0 1580.6817447447447u,0 1580.682744744745u,1.5 1581.6592847847846u,1.5 1581.6602847847848u,0 1582.6368248248248u,0 1582.637824824825u,1.5 1583.614364864865u,1.5 1583.6153648648651u,0 1584.5919049049048u,0 1584.592904904905u,1.5 1586.5469849849849u,1.5 1586.547984984985u,0 1587.524525025025u,0 1587.5255250250252u,1.5 1589.479605105105u,1.5 1589.4806051051053u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1603.1651656656657u,1.5 1603.1661656656659u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1607.0753258258258u,0 1607.076325825826u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1618.805806306306u,1.5 1618.8068063063063u,0 1619.7833463463462u,0 1619.7843463463464u,1.5 1621.7384264264263u,1.5 1621.7394264264265u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1650.0870875875873u,1.5 1650.0880875875876u,0 1651.0646276276275u,0 1651.0656276276277u,1.5 1652.0421676676676u,1.5 1652.0431676676678u,0 1662.795108108108u,0 1662.7961081081082u,1.5 1674.5255885885883u,1.5 1674.5265885885885u,0 1675.5031286286285u,0 1675.5041286286287u,1.5 1676.4806686686686u,1.5 1676.4816686686688u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1689.1886891891893u,1.5 1689.1896891891895u,0 1690.1662292292292u,0 1690.1672292292294u,1.5 1695.0539294294292u,1.5 1695.0549294294294u,0 1696.0314694694694u,0 1696.0324694694696u,1.5 1698.9640895895895u,1.5 1698.9650895895898u,0 1704.8293298298297u,0 1704.83032982983u,1.5 1705.8068698698698u,1.5 1705.80786986987u,0 1707.76194994995u,0 1707.76294994995u,1.5 1719.4924304304302u,1.5 1719.4934304304304u,0 1728.2902907907908u,0 1728.291290790791u,1.5 1729.2678308308307u,1.5 1729.268830830831u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1737.0881511511511u,1.5 1737.0891511511513u,0 1738.0656911911913u,0 1738.0666911911915u,1.5 1740.998311311311u,1.5 1740.9993113113112u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1752.7287917917918u,0 1752.729791791792u,1.5 1758.594032032032u,1.5 1758.5950320320321u,0 1759.571572072072u,0 1759.5725720720723u,1.5 1761.526652152152u,1.5 1761.5276521521523u,0 1767.3918923923923u,0 1767.3928923923925u,1.5 1768.3694324324322u,1.5 1768.3704324324324u,0 1771.3020525525524u,0 1771.3030525525526u,1.5 1781.0774529529529u,1.5 1781.078452952953u,0 1784.010073073073u,0 1784.0110730730732u,1.5 1784.987613113113u,1.5 1784.9886131131132u,0 1790.852853353353u,0 1790.8538533533533u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1794.7630135135132u,1.5 1794.7640135135134u,0 1795.7405535535534u,0 1795.7415535535536u,1.5 1802.5833338338336u,1.5 1802.5843338338339u,0 1803.5608738738738u,0 1803.561873873874u,1.5 1804.5384139139137u,1.5 1804.539413913914u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1823.1116746746745u,1.5 1823.1126746746747u,0 1824.0892147147147u,0 1824.0902147147149u,1.5 1826.0442947947947u,1.5 1826.045294794795u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1839.7298553553553u,0 1839.7308553553555u,1.5 1851.4603358358356u,1.5 1851.4613358358358u,0 1855.370495995996u,0 1855.3714959959962u,1.5 1856.3480360360359u,1.5 1856.349036036036u,0 1863.1908163163164u,0 1863.1918163163166u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1866.1234364364361u,0 1866.1244364364363u,1.5 1876.8763768768767u,1.5 1876.877376876877u,0 1877.853916916917u,0 1877.854916916917u,1.5 1878.8314569569568u,1.5 1878.832456956957u,0 1889.5843973973974u,0 1889.5853973973976u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1896.4271776776775u,0 1896.4281776776777u,1.5 1897.4047177177176u,1.5 1897.4057177177178u,0 1898.3822577577575u,0 1898.3832577577577u,1.5 1899.3597977977977u,1.5 1899.3607977977979u,0 1900.3373378378376u,0 1900.3383378378378u,1.5 1911.0902782782782u,1.5 1911.0912782782784u,0 1915.0004384384383u,0 1915.0014384384385u,1.5 1916.9555185185184u,1.5 1916.9565185185186u,0 1929.6635390390388u,0 1929.664539039039u,1.5 1930.641079079079u,1.5 1930.6420790790792u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1940.4164794794794u,1.5 1940.4174794794797u,0 1941.3940195195194u,0 1941.3950195195196u,1.5 1943.3490995995994u,1.5 1943.3500995995996u,0 1944.3266396396396u,0 1944.3276396396398u,1.5 1958.9897402402403u,1.5 1958.9907402402405u,0 1959.9672802802804u,0 1959.9682802802806u,1.5 1960.94482032032u,1.5 1960.9458203203203u,0 1961.9223603603602u,0 1961.9233603603604u,1.5 1964.8549804804804u,1.5 1964.8559804804806u,0 1965.8325205205203u,0 1965.8335205205206u,1.5 1967.7876006006004u,1.5 1967.7886006006006u,0 1968.7651406406405u,0 1968.7661406406407u,1.5 1970.7202207207204u,1.5 1970.7212207207206u,0 1971.6977607607605u,0 1971.6987607607607u,1.5 1974.630380880881u,1.5 1974.6313808808811u,0 1976.5854609609607u,0 1976.586460960961u,1.5 1977.5630010010009u,1.5 1977.564001001001u,0 1980.4956211211208u,0 1980.496621121121u,1.5 1981.473161161161u,1.5 1981.4741611611612u,0 1983.4282412412413u,0 1983.4292412412415u,1.5 1984.4057812812814u,1.5 1984.4067812812816u,0 1987.3384014014014u,0 1987.3394014014016u,1.5 1988.3159414414415u,1.5 1988.3169414414417u,0 1989.2934814814816u,0 1989.2944814814819u,1.5 1990.2710215215213u,1.5 1990.2720215215215u,0 1995.1587217217213u,0 1995.1597217217216u,1.5 1996.1362617617615u,1.5 1996.1372617617617u,0 1998.0913418418418u,0 1998.092341841842u,1.5 1999.068881881882u,1.5 1999.069881881882u,0 2007.8667422422423u,0 2007.8677422422425u,1.5 2008.8442822822824u,1.5 2008.8452822822826u,0 2014.7095225225223u,0 2014.7105225225225u,1.5 2015.6870625625625u,1.5 2015.6880625625627u,0 2021.5523028028026u,0 2021.5533028028028u,1.5 2022.5298428428428u,1.5 2022.530842842843u,0 2023.507382882883u,0 2023.508382882883u,1.5 2024.4849229229226u,1.5 2024.4859229229228u,0 2025.4624629629627u,0 2025.463462962963u,1.5 2026.4400030030029u,1.5 2026.441003003003u,0 2027.417543043043u,0 2027.4185430430432u,1.5 2028.3950830830831u,1.5 2028.3960830830833u,0 2029.3726231231228u,0 2029.373623123123u,1.5 2032.3052432432432u,1.5 2032.3062432432434u,0 2033.2827832832834u,0 2033.2837832832836u,1.5 2036.2154034034033u,1.5 2036.2164034034035u,0 2037.1929434434435u,0 2037.1939434434437u,1.5 2041.1031036036034u,1.5 2041.1041036036036u,0 2042.0806436436435u,0 2042.0816436436437u,1.5 2059.676364364364u,1.5 2059.677364364364u,0 2060.6539044044043u,0 2060.6549044044045u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2067.4966846846846u,1.5 2067.497684684685u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2070.429304804805u,1.5 2070.430304804805u,0 2086.0699454454452u,0 2086.0709454454454u,1.5 2091.9351856856856u,1.5 2091.936185685686u,0 2092.9127257257255u,0 2092.9137257257257u,1.5 2103.665666166166u,1.5 2103.666666166166u,0 2104.643206206206u,0 2104.644206206206u,1.5 2105.620746246246u,1.5 2105.6217462462464u,0 2120.2838468468467u,0 2120.284846846847u,1.5 2121.261386886887u,1.5 2121.2623868868873u,0 2123.216466966967u,0 2123.217466966967u,1.5 2134.946947447447u,1.5 2134.9479474474474u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2137.8795675675674u,1.5 2137.8805675675676u,0 2138.8571076076073u,0 2138.8581076076075u,1.5 2139.8346476476477u,1.5 2139.835647647648u,0 2149.610048048048u,0 2149.6110480480484u,1.5 2162.3180685685684u,1.5 2162.3190685685686u,0 2163.2956086086083u,0 2163.2966086086085u,1.5 2164.2731486486487u,1.5 2164.274148648649u,0 2174.048549049049u,0 2174.0495490490493u,1.5 2184.8014894894895u,1.5 2184.8024894894897u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2187.7341096096093u,1.5 2187.7351096096095u,0 2196.53196996997u,0 2196.53296996997u,1.5 2197.5095100100098u,1.5 2197.51051001001u,0 2198.48705005005u,0 2198.4880500500503u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2219.992930930931u,0 2219.993930930931u,1.5 2220.970470970971u,1.5 2220.971470970971u,0 2221.9480110110107u,0 2221.949011011011u,1.5 2227.813251251251u,1.5 2227.8142512512513u,0 2228.790791291291u,0 2228.7917912912912u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2230.745871371371u,0 2230.746871371371u,1.5 2231.7234114114112u,1.5 2231.7244114114114u,0 2238.5661916916915u,0 2238.5671916916917u,1.5 2239.543731731732u,1.5 2239.544731731732u,0 2240.5212717717714u,0 2240.5222717717716u,1.5 2241.4988118118117u,1.5 2241.499811811812u,0 2242.4763518518516u,0 2242.477351851852u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2254.2068323323324u,1.5 2254.2078323323326u,0 2260.0720725725723u,0 2260.0730725725725u,1.5 2268.869932932933u,1.5 2268.870932932933u,0 2269.847472972973u,0 2269.848472972973u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2280.600413413413u,0 2280.6014134134134u,1.5 2281.577953453453u,1.5 2281.5789534534533u,0 2282.5554934934935u,0 2282.5564934934937u,1.5 2290.3758138138137u,1.5 2290.376813813814u,0 2292.330893893894u,0 2292.331893893894u,1.5 2293.308433933934u,1.5 2293.309433933934u,0 2304.0613743743743u,0 2304.0623743743745u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2314.8143148148147u,0 2314.815314814815u,1.5 2316.769394894895u,1.5 2316.770394894895u,0 2317.746934934935u,0 2317.747934934935u,1.5 2318.724474974975u,1.5 2318.725474974975u,0 2324.589715215215u,0 2324.5907152152154u,1.5 2325.567255255255u,1.5 2325.5682552552553u,0 2327.5223353353354u,0 2327.5233353353356u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2340.2303558558556u,0 2340.231355855856u,1.5 2341.207895895896u,1.5 2341.208895895896u,0 2349.028216216216u,0 2349.0292162162164u,1.5 2350.005756256256u,1.5 2350.0067562562563u,0 2350.9832962962964u,0 2350.9842962962966u,1.5 2359.7811566566565u,1.5 2359.7821566566568u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2365.646396896897u,1.5 2365.647396896897u,0 2367.6014769769768u,0 2367.602476976977u,1.5 2368.5790170170167u,1.5 2368.580017017017u,0 2376.3993373373373u,0 2376.4003373373375u,1.5 2377.3768773773777u,1.5 2377.377877377378u,0 2380.3094974974974u,0 2380.3104974974976u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2397.905218218218u,1.5 2397.9062182182183u,0 2410.613238738739u,0 2410.614238738739u,1.5 2411.5907787787787u,1.5 2411.591778778779u,0 2412.5683188188186u,0 2412.569318818819u,1.5 2415.500938938939u,1.5 2415.501938938939u,0 2416.478478978979u,0 2416.4794789789794u,1.5 2432.119119619619u,1.5 2432.1201196196193u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2435.05173973974u,0 2435.05273973974u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.9843598598595u,0 2437.9853598598597u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2459.490240740741u,0 2459.491240740741u,1.5 2460.4677807807807u,1.5 2460.468780780781u,0 2461.4453208208206u,0 2461.446320820821u,1.5 2462.4228608608605u,1.5 2462.4238608608607u,0 2464.377940940941u,0 2464.378940940941u,1.5 2465.355480980981u,1.5 2465.3564809809814u,0 2466.3330210210206u,0 2466.334021021021u,1.5 2467.310561061061u,1.5 2467.311561061061u,0 2468.288101101101u,0 2468.289101101101u,1.5 2472.198261261261u,1.5 2472.199261261261u,0 2474.1533413413413u,0 2474.1543413413415u,1.5 2476.108421421421u,1.5 2476.1094214214213u,0 2478.0635015015014u,0 2478.0645015015016u,1.5 2482.9512017017014u,1.5 2482.9522017017016u,0 2483.9287417417418u,0 2483.929741741742u,1.5 2484.9062817817817u,1.5 2484.907281781782u,0 2485.8838218218216u,0 2485.884821821822u,1.5 2501.5244624624625u,1.5 2501.5254624624627u,0 2502.5020025025024u,0 2502.5030025025026u,1.5 2503.4795425425427u,1.5 2503.480542542543u,0 2504.4570825825826u,0 2504.458082582583u,1.5 2512.277402902903u,1.5 2512.278402902903u,0 2513.2549429429428u,0 2513.255942942943u,1.5 2517.165103103103u,1.5 2517.166103103103u,0 2518.1426431431432u,0 2518.1436431431434u,1.5 2519.120183183183u,1.5 2519.1211831831833u,0 2520.097723223223u,0 2520.0987232232233u,1.5 2522.0528033033033u,1.5 2522.0538033033035u,0 2523.0303433433432u,0 2523.0313433433435u,1.5 2524.985423423423u,1.5 2524.9864234234233u,0 2525.9629634634634u,0 2525.9639634634636u,1.5 2527.9180435435437u,1.5 2527.919043543544u,0 2528.8955835835836u,0 2528.896583583584u,1.5 2529.8731236236235u,1.5 2529.8741236236237u,0 2531.8282037037034u,0 2531.8292037037036u,1.5 2532.8057437437437u,1.5 2532.806743743744u,0 2533.7832837837836u,0 2533.784283783784u,1.5 2534.7608238238236u,1.5 2534.7618238238238u,0 2544.536224224224u,0 2544.5372242242242u,1.5 2545.513764264264u,1.5 2545.514764264264u,0 2554.3116246246245u,0 2554.3126246246247u,1.5 2555.2891646646644u,1.5 2555.2901646646646u,0 2558.2217847847846u,0 2558.222784784785u,1.5 2559.1993248248245u,1.5 2559.2003248248247u,0 2560.1768648648645u,0 2560.1778648648647u,1.5 2562.1319449449447u,1.5 2562.132944944945u,0 2565.064565065065u,0 2565.065565065065u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2567.019645145145u,0 2567.0206451451454u,1.5 2567.997185185185u,1.5 2567.9981851851853u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2586.5704459459457u,1.5 2586.571445945946u,0 2587.547985985986u,0 2587.5489859859863u,1.5 2588.5255260260255u,1.5 2588.5265260260257u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2608.0763268268265u,0 2608.0773268268267u,1.5 2619.8068073073073u,1.5 2619.8078073073075u,0 2620.784347347347u,0 2620.7853473473474u,1.5 2622.739427427427u,1.5 2622.740427427427u,0 2634.469907907908u,0 2634.470907907908u,1.5 2635.4474479479477u,1.5 2635.448447947948u,0 2637.402528028028u,0 2637.403528028028u,1.5 2650.1105485485486u,1.5 2650.111548548549u,0 2652.065628628629u,0 2652.066628628629u,1.5 2653.0431686686684u,1.5 2653.0441686686686u,0 2657.9308688688684u,0 2657.9318688688686u,1.5 2658.9084089089088u,1.5 2658.909408908909u,0 2659.8859489489487u,0 2659.886948948949u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2665.751189189189u,1.5 2665.7521891891893u,0 2666.7287292292294u,0 2666.7297292292296u,1.5 2672.5939694694694u,1.5 2672.5949694694696u,0 2673.5715095095093u,0 2673.5725095095095u,1.5 2674.5490495495496u,1.5 2674.55004954955u,0 2685.30198998999u,0 2685.3029899899902u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2689.21215015015u,1.5 2689.2131501501503u,0 2690.18969019019u,0 2690.1906901901903u,1.5 2694.09985035035u,1.5 2694.1008503503504u,0 2695.0773903903905u,0 2695.0783903903907u,1.5 2696.0549304304304u,1.5 2696.0559304304306u,0 2698.0100105105103u,0 2698.0110105105105u,1.5 2698.9875505505506u,1.5 2698.988550550551u,0 2699.9650905905905u,0 2699.9660905905907u,1.5 2700.942630630631u,1.5 2700.943630630631u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2710.718031031031u,1.5 2710.719031031031u,0 2711.695571071071u,0 2711.696571071071u,1.5 2718.538351351351u,1.5 2718.5393513513513u,0 2719.5158913913915u,0 2719.5168913913917u,1.5 2720.4934314314314u,1.5 2720.4944314314316u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2730.268831831832u,0 2730.269831831832u,1.5 2737.1116121121117u,1.5 2737.112612112112u,0 2738.089152152152u,0 2738.0901521521523u,1.5 2739.066692192192u,1.5 2739.067692192192u,0 2740.0442322322324u,0 2740.0452322322326u,1.5 2741.021772272272u,1.5 2741.022772272272u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2750.7971726726723u,0 2750.7981726726725u,1.5 2751.7747127127127u,1.5 2751.775712712713u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 2756.6624129129127u,1.5 2756.663412912913u,0 2757.6399529529526u,0 2757.640952952953u,1.5 2760.572573073073u,1.5 2760.573573073073u,0 2761.5501131131127u,0 2761.551113113113u,1.5 2762.527653153153u,1.5 2762.5286531531533u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2773.2805935935935u,0 2773.2815935935937u,1.5 2782.0784539539536u,1.5 2782.079453953954u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2801.6292547547546u,1.5 2801.630254754755u,0 2803.584334834835u,0 2803.585334834835u,1.5 2804.561874874875u,1.5 2804.562874874875u,0 2805.5394149149147u,0 2805.540414914915u,1.5 2806.5169549549546u,1.5 2806.517954954955u,0 2814.337275275275u,0 2814.338275275275u,1.5 2822.1575955955955u,1.5 2822.1585955955957u,0 2823.135135635636u,0 2823.136135635636u,1.5 2824.1126756756753u,1.5 2824.1136756756755u,0 2825.0902157157157u,0 2825.091215715716u,1.5 2826.0677557557556u,1.5 2826.068755755756u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2839.753316316316u,1.5 2839.7543163163164u,0 2840.730856356356u,0 2840.7318563563563u,1.5 2848.5511766766763u,1.5 2848.5521766766765u,0 2850.5062567567566u,0 2850.5072567567568u,1.5 2852.461336836837u,1.5 2852.462336836837u,0 2860.281657157157u,0 2860.2826571571572u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2865.169357357357u,1.5 2865.1703573573573u,0 2866.1468973973974u,0 2866.1478973973976u,1.5 2875.922297797798u,1.5 2875.923297797798u,0 2876.899837837838u,0 2876.900837837838u,1.5 2877.877377877878u,1.5 2877.8783778778784u,0 2878.8549179179176u,0 2878.855917917918u,1.5 2879.832457957958u,1.5 2879.833457957958u,0 2880.809997997998u,0 2880.810997997998u,1.5 2881.787538038038u,1.5 2881.788538038038u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2909.158659159159u,1.5 2909.159659159159u,0 2910.136199199199u,0 2910.137199199199u,1.5 2912.091279279279u,1.5 2912.0922792792794u,0 2913.068819319319u,0 2913.0698193193193u,1.5 2914.046359359359u,1.5 2914.0473593593592u,0 2930.66454004004u,0 2930.66554004004u,1.5 2931.64208008008u,1.5 2931.6430800800804u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2938.48486036036u,1.5 2938.48586036036u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2941.4174804804807u,0 2941.418480480481u,1.5 2942.39502052052u,1.5 2942.3960205205203u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 2958.035661161161u,1.5 2958.036661161161u,0 2959.013201201201u,0 2959.014201201201u,1.5 2962.923361361361u,1.5 2962.924361361361u,0 2963.9009014014014u,0 2963.9019014014016u,1.5 2965.8559814814816u,1.5 2965.856981481482u,0 2966.833521521521u,0 2966.8345215215213u,1.5 2968.7886016016014u,1.5 2968.7896016016016u,0 2969.7661416416418u,0 2969.767141641642u,1.5 2970.7436816816817u,1.5 2970.744681681682u,0 2971.7212217217216u,0 2971.722221721722u,1.5 2972.6987617617615u,1.5 2972.6997617617617u,0 2973.676301801802u,0 2973.677301801802u,1.5 2974.6538418418418u,1.5 2974.654841841842u,0 2979.541542042042u,0 2979.542542042042u,1.5 2980.519082082082u,1.5 2980.5200820820824u,0 2982.474162162162u,0 2982.475162162162u,1.5 2983.451702202202u,1.5 2983.452702202202u,0 2992.2495625625625u,0 2992.2505625625627u,1.5 2993.2271026026024u,1.5 2993.2281026026026u,0 3006.912663163163u,0 3006.913663163163u,1.5 3007.890203203203u,1.5 3007.891203203203u,0 3008.8677432432432u,0 3008.8687432432434u,1.5 3009.845283283283u,1.5 3009.8462832832834u,0 3010.822823323323u,0 3010.8238233233233u,1.5 3011.800363363363u,1.5 3011.801363363363u,0 3013.7554434434433u,0 3013.7564434434435u,1.5 3014.7329834834836u,1.5 3014.733983483484u,0 3016.6880635635634u,0 3016.6890635635636u,1.5 3017.6656036036034u,1.5 3017.6666036036036u,0 3018.6431436436437u,0 3018.644143643644u,1.5 3019.6206836836836u,1.5 3019.621683683684u,0 3022.553303803804u,0 3022.554303803804u,1.5 3024.508383883884u,1.5 3024.5093838838843u,0 3025.4859239239236u,0 3025.4869239239238u,1.5 3027.441004004004u,1.5 3027.442004004004u,0 3028.418544044044u,0 3028.4195440440444u,1.5 3029.396084084084u,1.5 3029.3970840840843u,0 3030.373624124124u,0 3030.3746241241242u,1.5 3032.328704204204u,1.5 3032.329704204204u,0 3033.306244244244u,0 3033.3072442442444u,1.5 3034.283784284284u,1.5 3034.2847842842843u,0 3035.261324324324u,0 3035.2623243243243u,1.5 3038.1939444444442u,1.5 3038.1949444444444u,0 3039.1714844844846u,0 3039.172484484485u,1.5 3042.1041046046043u,1.5 3042.1051046046045u,0 3043.0816446446447u,0 3043.082644644645u,1.5 3062.6324454454452u,1.5 3062.6334454454454u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3066.5426056056053u,0 3066.5436056056055u,1.5 3067.5201456456457u,1.5 3067.521145645646u,0 3084.138326326326u,0 3084.139326326326u,1.5 3085.115866366366u,1.5 3085.116866366366u,0 3088.0484864864866u,0 3088.049486486487u,1.5 3090.0035665665664u,1.5 3090.0045665665666u,0 3090.9811066066063u,0 3090.9821066066065u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3104.666667167167u,0 3104.667667167167u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3118.3522277277275u,0 3118.3532277277277u,1.5 3120.307307807808u,1.5 3120.308307807808u,0 3122.262387887888u,0 3122.2633878878883u,1.5 3125.195008008008u,1.5 3125.196008008008u,0 3126.172548048048u,0 3126.1735480480484u,1.5 3135.947948448448u,1.5 3135.9489484484484u,0 3147.678428928929u,0 3147.679428928929u,1.5 3148.655968968969u,1.5 3148.656968968969u,0 3151.588589089089u,0 3151.5895890890893u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3175.04955005005u,0 3175.0505500500503u,1.5 3177.0046301301304u,1.5 3177.0056301301306u,0 3177.98217017017u,0 3177.98317017017u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3196.555430930931u,0 3196.556430930931u,1.5 3197.532970970971u,1.5 3197.533970970971u,0 3198.5105110110107u,0 3198.511511011011u,1.5 3207.308371371371u,1.5 3207.309371371371u,0 3216.106231731732u,0 3216.107231731732u,1.5 3217.0837717717714u,1.5 3217.0847717717716u,0 3218.0613118118117u,0 3218.062311811812u,1.5 3219.0388518518516u,1.5 3219.039851851852u,0 3220.016391891892u,0 3220.017391891892u,1.5 3227.836712212212u,1.5 3227.8377122122124u,0 3228.814252252252u,0 3228.8152522522523u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3232.724412412412u,0 3232.7254124124124u,1.5 3233.701952452452u,1.5 3233.7029524524523u,0 3237.6121126126122u,0 3237.6131126126124u,1.5 3238.5896526526526u,1.5 3238.590652652653u,0 3239.5671926926925u,0 3239.5681926926927u,1.5 3240.544732732733u,1.5 3240.545732732733u,0 3241.5222727727723u,0 3241.5232727727725u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3259.1179934934935u,0 3259.1189934934937u,1.5 3260.0955335335334u,1.5 3260.0965335335336u,0 3262.050613613613u,0 3262.0516136136134u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3273.781094094094u,1.5 3273.782094094094u,0 3278.6687942942945u,0 3278.6697942942947u,1.5 3279.6463343343344u,1.5 3279.6473343343346u,0 3280.6238743743743u,0 3280.6248743743745u,1.5 3281.601414414414u,1.5 3281.6024144144144u,0 3283.5564944944945u,0 3283.5574944944947u,1.5 3290.3992747747743u,1.5 3290.4002747747745u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3294.309434934935u,1.5 3294.310434934935u,0 3302.129755255255u,0 3302.1307552552553u,1.5 3303.1072952952954u,1.5 3303.1082952952956u,0 3304.0848353353354u,0 3304.0858353353356u,1.5 3309.9500755755753u,1.5 3309.9510755755755u,0 3310.927615615615u,0 3310.9286156156154u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3325.590716216216u,0 3325.5917162162164u,1.5 3335.366116616616u,1.5 3335.3671166166164u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3349.0516771771768u,0 3349.052677177177u,1.5 3350.029217217217u,1.5 3350.0302172172173u,0 3351.006757257257u,0 3351.0077572572573u,1.5 3351.9842972972974u,1.5 3351.9852972972976u,0 3352.9618373373373u,0 3352.9628373373375u,1.5 3353.9393773773772u,1.5 3353.9403773773774u,0 3354.916917417417u,0 3354.9179174174174u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3365.6698578578576u,0 3365.6708578578578u,1.5 3366.647397897898u,1.5 3366.648397897898u,0 3378.3778783783787u,0 3378.378878378379u,1.5 3383.2655785785787u,1.5 3383.266578578579u,0 3384.243118618618u,0 3384.2441186186184u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3390.1083588588585u,0 3390.1093588588587u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.996059059059u,0 3394.997059059059u,1.5 3396.9511391391393u,1.5 3396.9521391391395u,0 3409.6591596596595u,0 3409.6601596596597u,1.5 3410.6366996996994u,1.5 3410.6376996996996u,0 3413.5693198198196u,0 3413.57031981982u,1.5 3415.5243998999u,1.5 3415.5253998999u,0 3417.47947997998u,0 3417.4804799799804u,1.5 3418.4570200200196u,1.5 3418.45802002002u,0 3419.43456006006u,0 3419.43556006006u,1.5 3431.1650405405403u,1.5 3431.1660405405405u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3434.0976606606605u,1.5 3434.0986606606607u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3436.052740740741u,1.5 3436.053740740741u,0 3455.6035415415413u,0 3455.6045415415415u,1.5 3456.5810815815817u,1.5 3456.582081581582u,0 3458.5361616616615u,0 3458.5371616616617u,1.5 3459.5137017017014u,1.5 3459.5147017017016u,0 3463.4238618618615u,0 3463.4248618618617u,1.5 3464.401401901902u,1.5 3464.402401901902u,0 3466.356481981982u,0 3466.3574819819823u,1.5 3468.311562062062u,1.5 3468.312562062062u,0 3469.289102102102u,0 3469.290102102102u,1.5 3471.244182182182u,1.5 3471.2451821821824u,0 3472.221722222222u,0 3472.2227222222223u,1.5 3475.1543423423423u,1.5 3475.1553423423425u,0 3476.1318823823826u,0 3476.132882382383u,1.5 3478.0869624624625u,1.5 3478.0879624624627u,0 3479.0645025025024u,0 3479.0655025025026u,1.5 3484.9297427427427u,1.5 3484.930742742743u,0 3485.9072827827827u,0 3485.908282782783u,1.5 3486.8848228228226u,1.5 3486.885822822823u,0 3487.8623628628625u,0 3487.8633628628627u,1.5 3488.839902902903u,1.5 3488.840902902903u,0 3489.8174429429428u,0 3489.818442942943u,1.5 3497.637763263263u,1.5 3497.638763263263u,0 3498.6153033033033u,0 3498.6163033033035u,1.5 3500.5703833833836u,1.5 3500.571383383384u,0 3501.547923423423u,0 3501.5489234234233u,1.5 3511.3233238238236u,1.5 3511.3243238238238u,0 3512.3008638638635u,0 3512.3018638638637u,1.5 3514.2559439439437u,1.5 3514.256943943944u,0 3515.233483983984u,0 3515.2344839839843u,1.5 3521.098724224224u,1.5 3521.0997242242242u,0 3522.076264264264u,0 3522.077264264264u,1.5 3524.0313443443442u,1.5 3524.0323443443444u,0 3525.986424424424u,0 3525.9874244244243u,1.5 3527.9415045045043u,1.5 3527.9425045045045u,0 3528.9190445445447u,0 3528.920044544545u,1.5 3529.8965845845846u,1.5 3529.897584584585u,0 3530.8741246246245u,0 3530.8751246246247u,1.5 3532.8292047047044u,1.5 3532.8302047047046u,0 3538.6944449449447u,0 3538.695444944945u,1.5 3539.671984984985u,1.5 3539.6729849849853u,0 3562.155405905906u,0 3562.156405905906u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.020646146146u,1.5 3568.0216461461464u,0 3568.998186186186u,0 3568.9991861861863u,1.5 3577.7960465465467u,1.5 3577.797046546547u,0 3578.7735865865866u,0 3578.774586586587u,1.5 3586.593906906907u,1.5 3586.594906906907u,0 3587.5714469469467u,0 3587.572446946947u,1.5 3588.548986986987u,1.5 3588.5499869869873u,0 3591.481607107107u,0 3591.482607107107u,1.5 3592.459147147147u,1.5 3592.4601471471474u,0 3603.2120875875876u,0 3603.213087587588u,1.5 3605.1671676676674u,1.5 3605.1681676676676u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3607.1222477477477u,1.5 3607.123247747748u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3621.785348348348u,1.5 3621.7863483483484u,0 3623.740428428428u,0 3623.741428428428u,1.5 3624.7179684684684u,1.5 3624.7189684684686u,0 3635.4709089089088u,0 3635.471908908909u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3637.425988988989u,0 3637.4269889889893u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3646.223849349349u,1.5 3646.2248493493494u,0 3647.2013893893895u,0 3647.2023893893897u,1.5 3651.1115495495496u,1.5 3651.11254954955u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3673.5949704704703u,1.5 3673.5959704704705u,0 3674.5725105105103u,0 3674.5735105105105u,1.5 3675.5500505505506u,1.5 3675.551050550551u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3688.258071071071u,0 3688.259071071071u,1.5 3697.0559314314314u,1.5 3697.0569314314316u,0 3699.9885515515516u,0 3699.989551551552u,1.5 3700.9660915915915u,1.5 3700.9670915915917u,0 3706.831331831832u,0 3706.832331831832u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3717.584272272272u,1.5 3717.585272272272u,0 3719.539352352352u,0 3719.5403523523523u,1.5 3720.5168923923925u,1.5 3720.5178923923927u,0 3721.4944324324324u,0 3721.4954324324326u,1.5 3722.4719724724723u,1.5 3722.4729724724725u,0 3730.292292792793u,0 3730.293292792793u,1.5 3732.2473728728723u,1.5 3732.2483728728726u,0 3733.2249129129127u,0 3733.225912912913u,1.5 3739.090153153153u,1.5 3739.0911531531533u,0 3740.067693193193u,0 3740.068693193193u,1.5 3741.0452332332334u,1.5 3741.0462332332336u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3757.6634139139137u,1.5 3757.664413913914u,0 3758.6409539539536u,0 3758.641953953954u,1.5 3759.618493993994u,1.5 3759.619493993994u,0 3760.596034034034u,0 3760.597034034034u,1.5 3761.573574074074u,1.5 3761.574574074074u,0 3772.326514514514u,0 3772.3275145145144u,1.5 3780.146834834835u,1.5 3780.147834834835u,0 3781.124374874875u,0 3781.125374874875u,1.5 3783.0794549549546u,1.5 3783.080454954955u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3802.6302557557556u,1.5 3802.631255755756u,0 3803.607795795796u,0 3803.608795795796u,1.5 3804.585335835836u,1.5 3804.586335835836u,0 3806.5404159159157u,0 3806.541415915916u,1.5 3807.5179559559556u,1.5 3807.518955955956u,0 3812.405656156156u,0 3812.4066561561563u,1.5 3813.383196196196u,1.5 3813.384196196196u,0 3814.3607362362363u,0 3814.3617362362365u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3816.315816316316u,0 3816.3168163163164u,1.5 3817.293356356356u,1.5 3817.2943563563563u,0 3818.2708963963964u,0 3818.2718963963966u,1.5 3825.1136766766763u,1.5 3825.1146766766765u,0 3826.0912167167166u,0 3826.092216716717u,1.5 3827.0687567567566u,1.5 3827.0697567567568u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3836.844157157157u,1.5 3836.8451571571572u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 3847.5970975975974u,1.5 3847.5980975975976u,0 3848.574637637638u,0 3848.575637637638u,1.5 3850.5297177177176u,1.5 3850.530717717718u,0 3851.5072577577575u,0 3851.5082577577577u,1.5 3852.484797797798u,1.5 3852.485797797798u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3876.923298798799u,1.5 3876.924298798799u,0 3877.900838838839u,0 3877.901838838839u,1.5 3879.8559189189186u,1.5 3879.856918918919u,0 3887.6762392392393u,0 3887.6772392392395u,1.5 3888.653779279279u,1.5 3888.6547792792794u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3895.4965595595595u,0 3895.4975595595597u,1.5 3913.09228028028u,1.5 3913.0932802802804u,0 3914.06982032032u,0 3914.0708203203203u,1.5 3915.0473603603605u,1.5 3915.0483603603607u,0 3917.00244044044u,0 3917.00344044044u,1.5 3917.9799804804807u,1.5 3917.980980480481u,0 3933.6206211211206u,0 3933.621621121121u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3938.508321321321u,1.5 3938.5093213213213u,0 3939.4858613613615u,0 3939.4868613613617u,1.5 3960.991742242242u,1.5 3960.992742242242u,0 3961.969282282282u,0 3961.9702822822824u,1.5 3962.946822322322u,1.5 3962.9478223223223u,0 3963.9243623623624u,0 3963.9253623623626u,1.5 3965.879442442442u,1.5 3965.880442442442u,0 3966.8569824824826u,0 3966.857982482483u,1.5 3967.834522522522u,1.5 3967.8355225225223u,0 3969.7896026026024u,0 3969.7906026026026u,1.5 3972.7222227227226u,1.5 3972.7232227227228u,0 3973.699762762763u,0 3973.700762762763u,1.5 3974.677302802803u,1.5 3974.678302802803u,0 3975.6548428428423u,0 3975.6558428428425u,1.5 3977.6099229229226u,1.5 3977.610922922923u,0 3980.5425430430428u,0 3980.543543043043u,1.5 3981.520083083083u,1.5 3981.5210830830833u,0 3982.4976231231226u,0 3982.498623123123u,1.5 3983.4751631631634u,1.5 3983.4761631631636u,0 3989.3404034034033u,0 3989.3414034034035u,1.5 3990.317943443443u,1.5 3990.318943443443u,0 3998.138263763764u,0 3998.139263763764u,1.5 3999.115803803804u,1.5 3999.116803803804u,0 4013.7789044044043u,0 4013.7799044044045u,1.5 4014.756444444444u,1.5 4014.757444444444u,0 4016.711524524524u,0 4016.7125245245243u,1.5 4017.689064564565u,1.5 4017.690064564565u,0 4020.6216846846846u,0 4020.622684684685u,1.5 4021.5992247247245u,1.5 4021.6002247247247u,0 4024.5318448448443u,0 4024.5328448448445u,1.5 4026.4869249249246u,1.5 4026.4879249249248u,0 4027.4644649649654u,0 4027.4654649649656u,1.5 4028.442005005005u,1.5 4028.443005005005u,0 4029.4195450450447u,0 4029.420545045045u,1.5 4030.397085085085u,1.5 4030.3980850850853u,0 4031.374625125125u,0 4031.375625125125u,1.5 4033.329705205205u,1.5 4033.330705205205u,0 4035.284785285285u,0 4035.2857852852853u,1.5 4037.2398653653654u,1.5 4037.2408653653656u,0 4038.2174054054053u,0 4038.2184054054055u,1.5 4039.194945445445u,1.5 4039.195945445445u,0 4040.1724854854856u,0 4040.173485485486u,1.5 4043.1051056056053u,1.5 4043.1061056056055u,0 4044.0826456456452u,0 4044.0836456456454u,1.5 4057.768206206206u,1.5 4057.769206206206u,0 4058.7457462462457u,0 4058.746746246246u,1.5 4061.6783663663664u,1.5 4061.6793663663666u,0 4062.6559064064063u,0 4062.6569064064065u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4065.588526526526u,0 4065.5895265265262u,1.5 4066.566066566567u,1.5 4066.567066566567u,0 4067.5436066066063u,0 4067.5446066066065u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4080.251627127127u,0 4080.252627127127u,1.5 4081.2291671671674u,1.5 4081.2301671671676u,0 4084.161787287287u,0 4084.1627872872873u,1.5 4085.139327327327u,1.5 4085.140327327327u,0 4086.1168673673674u,0 4086.1178673673676u,1.5 4087.0944074074073u,1.5 4087.0954074074075u,0 4089.0494874874876u,0 4089.0504874874878u,1.5 4093.9371876876876u,1.5 4093.938187687688u,0 4094.9147277277275u,0 4094.9157277277277u,1.5 4101.757508008008u,1.5 4101.758508008008u,0 4102.735048048047u,0 4102.736048048047u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4105.667668168168u,0 4105.668668168169u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4119.353228728728u,0 4119.354228728728u,1.5 4120.330768768769u,1.5 4120.3317687687695u,0 4122.285848848848u,0 4122.286848848848u,1.5 4124.240928928929u,1.5 4124.241928928929u,0 4125.218468968969u,0 4125.2194689689695u,1.5 4134.993869369369u,1.5 4134.99486936937u,0 4137.9264894894895u,0 4137.92748948949u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4146.724349849849u,0 4146.725349849849u,1.5 4147.70188988989u,1.5 4147.70288988989u,0 4148.67942992993u,0 4148.68042992993u,1.5 4149.65696996997u,1.5 4149.6579699699705u,0 4150.63451001001u,0 4150.63551001001u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4172.140390890891u,0 4172.141390890891u,1.5 4173.117930930931u,1.5 4173.118930930931u,0 4174.095470970971u,0 4174.0964709709715u,1.5 4183.870871371371u,1.5 4183.8718713713715u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4193.646271771772u,0 4193.6472717717725u,1.5 4194.623811811812u,1.5 4194.624811811812u,0 4197.556431931932u,0 4197.557431931932u,1.5 4198.533971971972u,1.5 4198.5349719719725u,0 4199.511512012012u,0 4199.512512012012u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4209.286912412412u,1.5 4209.287912412412u,0 4219.062312812813u,0 4219.063312812813u,1.5 4225.9050930930935u,1.5 4225.906093093094u,0 4226.882633133133u,0 4226.883633133133u,1.5 4229.815253253253u,1.5 4229.816253253253u,0 4236.658033533533u,0 4236.659033533533u,1.5 4237.635573573573u,1.5 4237.6365735735735u,0 4238.613113613614u,0 4238.614113613614u,1.5 4239.590653653653u,1.5 4239.591653653653u,0 4240.5681936936935u,0 4240.569193693694u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4260.1189944944945u,0 4260.119994494495u,1.5 4261.096534534534u,1.5 4261.097534534534u,0 4262.074074574574u,0 4262.0750745745745u,1.5 4268.916854854855u,1.5 4268.917854854855u,0 4270.871934934935u,0 4270.872934934935u,1.5 4272.827015015015u,1.5 4272.828015015015u,0 4282.602415415415u,0 4282.603415415415u,1.5 4289.4451956956955u,1.5 4289.446195695696u,0 4290.422735735735u,0 4290.423735735735u,1.5 4292.377815815816u,1.5 4292.378815815816u,0 4293.355355855856u,0 4293.356355855856u,1.5 4294.3328958958955u,1.5 4294.333895895896u,0 4303.130756256257u,0 4303.131756256257u,1.5 4313.8836966966965u,1.5 4313.884696696697u,0 4322.681557057057u,0 4322.682557057057u,1.5 4323.659097097097u,1.5 4323.660097097098u,0 4326.591717217217u,0 4326.592717217217u,1.5 4327.569257257258u,1.5 4327.570257257258u,0 4328.546797297297u,0 4328.547797297298u,1.5 4336.367117617618u,1.5 4336.368117617618u,0 4337.344657657658u,0 4337.345657657658u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4342.232357857858u,1.5 4342.233357857858u,0 4347.120058058058u,0 4347.121058058058u,1.5 4348.097598098098u,1.5 4348.098598098099u,0 4351.030218218218u,0 4351.031218218218u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4362.760698698698u,0 4362.761698698699u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4368.625938938939u,0 4368.626938938939u,1.5 4369.603478978979u,1.5 4369.604478978979u,0 4373.513639139139u,0 4373.514639139139u,1.5 4374.491179179179u,1.5 4374.492179179179u,0 4376.44625925926u,0 4376.44725925926u,1.5 4377.423799299299u,1.5 4377.4247992993u,0 4379.378879379379u,0 4379.379879379379u,1.5 4390.13181981982u,1.5 4390.13281981982u,0 4391.10935985986u,0 4391.11035985986u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.99706006006u,1.5 4395.99806006006u,0 4411.6377007007u,0 4411.638700700701u,1.5 4412.61524074074u,1.5 4412.61624074074u,0 4414.570320820821u,0 4414.571320820821u,1.5 4416.5254009009u,1.5 4416.526400900901u,0 4417.502940940941u,0 4417.503940940941u,1.5 4418.480480980981u,1.5 4418.481480980981u,0 4419.458021021021u,0 4419.459021021021u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4438.031281781782u,1.5 4438.032281781782u,0 4440.963901901901u,0 4440.964901901902u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4456.604542542542u,0 4456.605542542542u,1.5 4457.582082582582u,1.5 4457.583082582582u,0 4462.469782782783u,0 4462.470782782783u,1.5 4463.447322822823u,1.5 4463.448322822823u,0 4465.402402902902u,0 4465.403402902903u,1.5 4466.379942942943u,1.5 4466.380942942943u,0 4467.357482982983u,0 4467.358482982983u,1.5 4468.335023023023u,1.5 4468.336023023023u,0 4469.312563063063u,0 4469.313563063063u,1.5 4470.290103103103u,1.5 4470.2911031031035u,0 4471.267643143143u,0 4471.268643143143u,1.5 4472.245183183183u,1.5 4472.246183183183u,0 4473.222723223223u,0 4473.223723223223u,1.5 4476.155343343343u,1.5 4476.156343343343u,0 4478.1104234234235u,0 4478.111423423424u,1.5 4479.087963463464u,1.5 4479.088963463464u,0 4480.065503503503u,0 4480.066503503504u,1.5 4488.863363863864u,1.5 4488.864363863864u,0 4489.840903903903u,0 4489.841903903904u,1.5 4490.818443943944u,1.5 4490.819443943944u,0 4491.795983983984u,0 4491.796983983984u,1.5 4492.773524024024u,1.5 4492.774524024024u,0 4493.751064064064u,0 4493.752064064064u,1.5 4494.728604104104u,1.5 4494.7296041041045u,0 4495.706144144144u,0 4495.707144144144u,1.5 4502.5489244244245u,1.5 4502.549924424425u,0 4503.526464464465u,0 4503.527464464465u,1.5 4505.481544544544u,1.5 4505.482544544544u,0 4506.459084584585u,0 4506.460084584585u,1.5 4516.234484984985u,1.5 4516.235484984985u,0 4517.212025025025u,0 4517.213025025025u,1.5 4519.167105105105u,1.5 4519.1681051051055u,0 4520.144645145145u,0 4520.145645145145u,1.5 4521.122185185185u,1.5 4521.123185185185u,0 4523.077265265266u,0 4523.078265265266u,1.5 4524.054805305305u,1.5 4524.0558053053055u,0 4525.032345345345u,0 4525.033345345345u,1.5 4526.009885385385u,1.5 4526.010885385385u,0 4526.9874254254255u,0 4526.988425425426u,1.5 4528.942505505505u,1.5 4528.9435055055055u,0 4530.897585585586u,0 4530.898585585586u,1.5 4532.852665665666u,1.5 4532.853665665666u,0 4534.807745745745u,0 4534.808745745745u,1.5 4535.785285785786u,1.5 4535.786285785786u,0 4565.111486986987u,0 4565.112486986987u,1.5 4566.0890270270265u,1.5 4566.090027027027u,0 4567.066567067067u,0 4567.067567067067u,1.5 4584.662287787788u,1.5 4584.663287787788u,0 4585.6398278278275u,0 4585.640827827828u,1.5 4586.617367867868u,1.5 4586.618367867868u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4609.100788788789u,1.5 4609.101788788789u,0 4610.0783288288285u,0 4610.079328828829u,1.5 4620.83126926927u,1.5 4620.83226926927u,0 4623.763889389389u,0 4623.764889389389u,1.5 4624.741429429429u,1.5 4624.74242942943u,0 4635.49436986987u,0 4635.49536986987u,1.5 4636.471909909909u,1.5 4636.4729099099095u,0 4637.44944994995u,0 4637.45044994995u,1.5 4648.20239039039u,1.5 4648.20339039039u,0 4649.17993043043u,0 4649.180930430431u,1.5 4651.13501051051u,1.5 4651.1360105105105u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4675.573511511511u,1.5 4675.574511511511u,0 4686.326451951952u,0 4686.327451951952u,1.5 4696.101852352352u,1.5 4696.102852352352u,0 4698.056932432432u,0 4698.057932432433u,1.5 4699.034472472473u,1.5 4699.035472472473u,0 4700.989552552552u,0 4700.990552552552u,1.5 4701.967092592593u,1.5 4701.968092592593u,0 4704.899712712712u,0 4704.900712712712u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4715.652653153153u,1.5 4715.653653153153u,0 4716.630193193193u,0 4716.631193193193u,1.5 4718.585273273274u,1.5 4718.586273273274u,0 4719.562813313313u,0 4719.563813313313u,1.5 4720.540353353353u,1.5 4720.541353353353u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4731.293293793794u,1.5 4731.294293793794u,0 4732.270833833833u,0 4732.271833833834u,1.5 4739.113614114114u,1.5 4739.114614114114u,0 4740.091154154154u,0 4740.092154154154u,1.5 4741.068694194194u,1.5 4741.069694194194u,0 4742.046234234233u,0 4742.047234234234u,1.5 4743.023774274275u,1.5 4743.024774274275u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4759.6419549549555u,1.5 4759.642954954956u,0 4760.619494994995u,0 4760.620494994995u,1.5 4761.597035035034u,1.5 4761.598035035035u,0 4768.439815315315u,0 4768.440815315315u,1.5 4769.4173553553555u,1.5 4769.418355355356u,0 4771.372435435435u,0 4771.373435435436u,1.5 4782.125375875876u,1.5 4782.126375875876u,0 4783.102915915916u,0 4783.103915915916u,1.5 4784.0804559559565u,1.5 4784.081455955957u,0 4793.8558563563565u,0 4793.856856356357u,1.5 4802.653716716716u,1.5 4802.654716716716u,0 4803.6312567567575u,0 4803.632256756758u,1.5 4805.586336836836u,1.5 4805.587336836837u,0 4806.563876876877u,0 4806.564876876877u,1.5 4807.541416916917u,1.5 4807.542416916917u,0 4815.361737237236u,0 4815.362737237237u,1.5 4825.137137637637u,1.5 4825.138137637638u,0 4826.114677677678u,0 4826.115677677678u,1.5 4828.069757757758u,1.5 4828.070757757759u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4840.777778278279u,1.5 4840.778778278279u,0 4841.755318318318u,0 4841.756318318318u,1.5 4848.598098598599u,1.5 4848.599098598599u,0 4849.575638638638u,0 4849.5766386386385u,1.5 4852.508258758759u,1.5 4852.50925875876u,0 4863.261199199199u,0 4863.262199199199u,1.5 4864.238739239238u,1.5 4864.239739239239u,0 4866.193819319319u,0 4866.194819319319u,1.5 4875.969219719719u,1.5 4875.970219719719u,0 4876.94675975976u,0 4876.947759759761u,1.5 4877.9242997998u,1.5 4877.9252997998u,0 4878.901839839839u,0 4878.9028398398395u,1.5 4879.87937987988u,1.5 4879.88037987988u,0 4880.85691991992u,0 4880.85791991992u,1.5 4881.83445995996u,1.5 4881.835459959961u,0 4891.6098603603605u,0 4891.610860360361u,1.5 4892.5874004004u,1.5 4892.5884004004u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4894.542480480481u,1.5 4894.543480480481u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4898.45264064064u,1.5 4898.4536406406405u,0 4899.430180680681u,0 4899.431180680681u,1.5 4912.138201201201u,1.5 4912.139201201201u,0 4913.11574124124u,0 4913.116741241241u,1.5 4914.093281281282u,1.5 4914.094281281282u,0 4915.070821321321u,0 4915.071821321321u,1.5 4916.0483613613615u,1.5 4916.049361361362u,0 4917.025901401401u,0 4917.026901401401u,1.5 4918.003441441441u,1.5 4918.0044414414415u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4938.531782282283u,0 4938.532782282283u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 4941.464402402402u,0 4941.465402402402u,1.5 4965.902903403403u,1.5 4965.903903403403u,0 4966.880443443443u,0 4966.8814434434435u,1.5 4968.835523523523u,1.5 4968.836523523523u,0 4970.790603603604u,0 4970.791603603604u,1.5 4971.768143643643u,1.5 4971.7691436436435u,0 4972.745683683684u,0 4972.746683683684u,1.5 4973.723223723723u,1.5 4973.724223723723u,0 4974.700763763764u,0 4974.701763763765u,1.5 4975.678303803804u,1.5 4975.679303803804u,0 4976.655843843843u,0 4976.6568438438435u,1.5 4977.633383883884u,1.5 4977.634383883884u,0 4979.588463963964u,0 4979.589463963965u,1.5 4980.566004004004u,1.5 4980.567004004004u,0 4983.498624124124u,0 4983.499624124124u,1.5 4984.476164164164u,1.5 4984.477164164165u,0 4986.431244244243u,0 4986.4322442442435u,1.5 4987.408784284285u,1.5 4987.409784284285u,0 4989.363864364364u,0 4989.364864364365u,1.5 4990.341404404404u,1.5 4990.342404404404u,0 4992.296484484485u,0 4992.297484484485u,1.5 4993.274024524524u,1.5 4993.275024524524u,0 4996.206644644644u,0 4996.2076446446445u,1.5 4997.184184684685u,1.5 4997.185184684685u,0 5007.937125125125u,0 5007.938125125125u,1.5 5008.914665165165u,1.5 5008.915665165166u,0 5014.779905405405u,0 5014.780905405405u,1.5 5015.757445445445u,1.5 5015.758445445445u,0 5016.734985485486u,0 5016.735985485486u,1.5 5017.712525525525u,1.5 5017.713525525525u,0 5021.622685685686u,0 5021.623685685686u,1.5 5022.600225725725u,1.5 5022.601225725725u,0 5024.555305805806u,0 5024.556305805806u,1.5 5025.532845845845u,1.5 5025.5338458458455u,0 5027.487925925926u,0 5027.488925925926u,1.5 5028.465465965966u,1.5 5028.466465965967u,0 5029.443006006006u,0 5029.444006006006u,1.5 5030.420546046045u,1.5 5030.4215460460455u,0 5031.398086086087u,0 5031.399086086087u,1.5 5033.353166166166u,1.5 5033.354166166167u,0 5035.308246246245u,0 5035.3092462462455u,1.5 5057.791667167167u,1.5 5057.792667167168u,0 5058.769207207207u,0 5058.770207207207u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5064.634447447447u,1.5 5064.635447447447u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5086.140328328328u,0 5086.141328328328u,1.5 5087.117868368368u,1.5 5087.118868368369u,0 5088.095408408408u,0 5088.096408408408u,1.5 5090.050488488489u,1.5 5090.051488488489u,0 5092.005568568568u,0 5092.006568568569u,1.5 5092.983108608609u,1.5 5092.984108608609u,0 5093.960648648648u,0 5093.961648648648u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5120.354229729729u,0 5120.355229729729u,1.5 5121.33176976977u,1.5 5121.3327697697705u,0 5123.286849849849u,0 5123.287849849849u,1.5 5124.26438988989u,1.5 5124.26538988989u,0 5125.24192992993u,0 5125.24292992993u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5135.99487037037u,0 5135.9958703703705u,1.5 5136.97241041041u,1.5 5136.97341041041u,0 5149.680430930931u,0 5149.681430930931u,1.5 5150.657970970971u,1.5 5150.6589709709715u,0 5152.61305105105u,0 5152.61405105105u,1.5 5160.433371371371u,1.5 5160.4343713713715u,0 5161.410911411411u,0 5161.411911411411u,1.5 5162.388451451451u,1.5 5162.389451451451u,0 5171.186311811812u,0 5171.187311811812u,1.5 5172.163851851851u,1.5 5172.164851851851u,0 5174.118931931932u,0 5174.119931931932u,1.5 5176.074012012012u,1.5 5176.075012012012u,0 5177.051552052051u,0 5177.052552052051u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5194.647272772773u,0 5194.648272772773u,1.5 5195.624812812813u,1.5 5195.625812812813u,0 5198.557432932933u,0 5198.558432932933u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5218.108233733733u,0 5218.109233733733u,1.5 5220.063313813814u,1.5 5220.064313813814u,0 5221.040853853853u,0 5221.041853853853u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5232.771334334334u,1.5 5232.772334334334u,0 5237.659034534534u,0 5237.660034534534u,1.5 5238.636574574574u,1.5 5238.6375745745745u,0 5240.591654654654u,0 5240.592654654654u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5258.187375375375u,0 5258.1883753753755u,1.5 5259.164915415415u,1.5 5259.165915415415u,0 5260.142455455456u,0 5260.143455455456u,1.5 5261.1199954954955u,1.5 5261.120995495496u,0 5262.097535535535u,0 5262.098535535535u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5280.670796296296u,0 5280.671796296297u,1.5 5281.648336336336u,1.5 5281.649336336336u,0 5282.625876376376u,0 5282.6268763763765u,1.5 5283.603416416417u,1.5 5283.604416416417u,0 5284.580956456457u,0 5284.581956456457u,1.5 5289.468656656657u,1.5 5289.469656656657u,0 5290.4461966966965u,0 5290.447196696697u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5294.356356856857u,0 5294.357356856857u,1.5 5295.3338968968965u,1.5 5295.334896896897u,0 5299.244057057057u,0 5299.245057057057u,1.5 5300.221597097097u,1.5 5300.222597097098u,0 5302.176677177177u,0 5302.177677177177u,1.5 5303.154217217217u,1.5 5303.155217217217u,0 5304.131757257258u,0 5304.132757257258u,1.5 5305.109297297297u,1.5 5305.110297297298u,0 5306.086837337337u,0 5306.087837337337u,1.5 5312.929617617618u,1.5 5312.930617617618u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5326.615178178178u,0 5326.616178178178u,1.5 5327.592718218218u,1.5 5327.593718218218u,0 5328.570258258259u,0 5328.571258258259u,1.5 5337.368118618619u,1.5 5337.369118618619u,0 5338.345658658659u,0 5338.346658658659u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5351.053679179179u,0 5351.054679179179u,1.5 5352.031219219219u,1.5 5352.032219219219u,0 5353.00875925926u,0 5353.00975925926u,1.5 5354.963839339339u,1.5 5354.964839339339u,0 5355.941379379379u,0 5355.942379379379u,1.5 5362.78415965966u,1.5 5362.78515965966u,0 5363.761699699699u,0 5363.7626996997u,1.5 5364.739239739739u,1.5 5364.740239739739u,0 5366.69431981982u,0 5366.69531981982u,1.5 5367.67185985986u,1.5 5367.67285985986u,0 5376.46972022022u,0 5376.47072022022u,1.5 5377.447260260261u,1.5 5377.448260260261u,0 5378.4248003003u,0 5378.425800300301u,1.5 5394.065440940941u,1.5 5394.066440940941u,0 5395.042980980981u,0 5395.043980980981u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5396.998061061061u,0 5396.999061061061u,1.5 5397.975601101101u,1.5 5397.976601101102u,0 5398.953141141141u,0 5398.954141141141u,1.5 5399.930681181181u,1.5 5399.931681181181u,0 5407.751001501501u,0 5407.752001501502u,1.5 5408.728541541541u,1.5 5408.729541541541u,0 5410.683621621622u,0 5410.684621621622u,1.5 5411.661161661662u,1.5 5411.662161661662u,0 5413.616241741741u,0 5413.617241741741u,1.5 5430.2344224224225u,1.5 5430.235422422423u,0 5431.211962462463u,0 5431.212962462463u,1.5 5432.189502502502u,1.5 5432.190502502503u,0 5433.167042542542u,0 5433.168042542542u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5438.054742742742u,0 5438.055742742742u,1.5 5439.032282782783u,1.5 5439.033282782783u,0 5440.009822822823u,0 5440.010822822823u,1.5 5440.987362862863u,1.5 5440.988362862863u,0 5444.897523023023u,0 5444.898523023023u,1.5 5445.875063063063u,1.5 5445.876063063063u,0 5461.515703703703u,0 5461.516703703704u,1.5 5462.493243743743u,1.5 5462.494243743743u,0 5464.448323823824u,0 5464.449323823824u,1.5 5465.425863863864u,1.5 5465.426863863864u,0 5470.313564064064u,0 5470.314564064064u,1.5 5471.291104104104u,1.5 5471.2921041041045u,0 5473.246184184184u,0 5473.247184184184u,1.5 5474.223724224224u,1.5 5474.224724224224u,0 5475.201264264265u,0 5475.202264264265u,1.5 5478.133884384384u,1.5 5478.134884384384u,0 5479.1114244244245u,0 5479.112424424425u,1.5 5481.066504504504u,1.5 5481.0675045045045u,0 5482.044044544544u,0 5482.045044544544u,1.5 5483.021584584585u,1.5 5483.022584584585u,0 5483.9991246246245u,0 5484.000124624625u,1.5 5484.976664664665u,1.5 5484.977664664665u,0 5485.954204704704u,0 5485.955204704705u,1.5 5488.8868248248245u,1.5 5488.887824824825u,0 5489.864364864865u,0 5489.865364864865u,1.5 5492.796984984985u,1.5 5492.797984984985u,0 5493.774525025025u,0 5493.775525025025u,1.5 5495.729605105105u,1.5 5495.7306051051055u,0 5496.707145145145u,0 5496.708145145145u,1.5 5499.639765265266u,1.5 5499.640765265266u,0 5500.617305305305u,0 5500.6183053053055u,1.5 5510.392705705705u,1.5 5510.3937057057055u,0 5511.370245745745u,0 5511.371245745745u,1.5 5515.280405905905u,1.5 5515.281405905906u,0 5516.257945945946u,0 5516.258945945946u,1.5 5517.235485985986u,1.5 5517.236485985986u,0 5518.213026026026u,0 5518.214026026026u,1.5 5520.168106106106u,1.5 5520.1691061061065u,0 5521.145646146146u,0 5521.146646146146u,1.5 5524.078266266267u,1.5 5524.079266266267u,0 5525.055806306306u,0 5525.0568063063065u,1.5 5526.033346346346u,1.5 5526.034346346346u,0 5527.010886386386u,0 5527.011886386386u,1.5 5527.9884264264265u,1.5 5527.989426426427u,0 5529.943506506506u,0 5529.9445065065065u,1.5 5530.921046546546u,1.5 5530.922046546546u,0 5531.898586586587u,0 5531.899586586587u,1.5 5533.853666666667u,1.5 5533.854666666667u,0 5540.696446946947u,0 5540.697446946947u,1.5 5541.673986986987u,1.5 5541.674986986987u,0 5558.292167667668u,0 5558.293167667668u,1.5 5559.269707707707u,1.5 5559.2707077077075u,0 5562.2023278278275u,0 5562.203327827828u,1.5 5563.179867867868u,1.5 5563.180867867868u,0 5566.112487987988u,0 5566.113487987988u,1.5 5567.0900280280275u,1.5 5567.091028028028u,0 5568.067568068068u,0 5568.068568068068u,1.5 5570.022648148148u,1.5 5570.023648148148u,0 5571.000188188188u,0 5571.001188188188u,1.5 5584.685748748749u,1.5 5584.686748748749u,0 5585.663288788789u,0 5585.664288788789u,1.5 5586.6408288288285u,1.5 5586.641828828829u,0 5587.618368868869u,0 5587.619368868869u,1.5 5589.573448948949u,1.5 5589.574448948949u,0 5600.326389389389u,0 5600.327389389389u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5605.21408958959u,0 5605.21508958959u,1.5 5608.146709709709u,1.5 5608.1477097097095u,0 5609.12424974975u,0 5609.12524974975u,1.5 5620.8547302302295u,1.5 5620.85573023023u,0 5621.832270270271u,0 5621.833270270271u,1.5 5623.78735035035u,1.5 5623.78835035035u,0 5633.562750750751u,0 5633.563750750751u,1.5 5634.540290790791u,1.5 5634.541290790791u,0 5636.495370870871u,0 5636.496370870871u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5638.450450950951u,0 5638.451450950951u,1.5 5648.225851351351u,1.5 5648.226851351351u,0 5649.203391391391u,0 5649.204391391391u,1.5 5650.180931431431u,1.5 5650.181931431432u,0 5651.158471471472u,0 5651.159471471472u,1.5 5652.136011511511u,1.5 5652.137011511511u,0 5653.113551551551u,0 5653.114551551551u,1.5 5654.091091591592u,1.5 5654.092091591592u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5664.8440320320315u,1.5 5664.845032032032u,0 5665.821572072072u,0 5665.822572072072u,1.5 5675.596972472473u,1.5 5675.597972472473u,0 5676.574512512512u,0 5676.575512512512u,1.5 5677.552052552552u,1.5 5677.553052552552u,0 5682.439752752753u,0 5682.440752752753u,1.5 5683.417292792793u,1.5 5683.418292792793u,0 5685.372372872873u,0 5685.373372872873u,1.5 5688.304992992993u,1.5 5688.305992992993u,0 5689.282533033032u,0 5689.283533033033u,1.5 5695.147773273274u,1.5 5695.148773273274u,0 5696.125313313313u,0 5696.126313313313u,1.5 5699.057933433433u,1.5 5699.058933433434u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5715.676114114114u,1.5 5715.677114114114u,0 5716.653654154154u,0 5716.654654154154u,1.5 5718.608734234233u,1.5 5718.609734234234u,0 5727.406594594595u,0 5727.407594594595u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5740.114615115115u,1.5 5740.115615115115u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 5758.687875875876u,1.5 5758.688875875876u,0 5759.665415915916u,0 5759.666415915916u,1.5 5760.6429559559565u,1.5 5760.643955955957u,0 5761.620495995996u,0 5761.621495995996u,1.5 5762.598036036035u,1.5 5762.599036036036u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5772.373436436436u,0 5772.374436436437u,1.5 5778.238676676677u,1.5 5778.239676676677u,0 5779.216216716716u,0 5779.217216716716u,1.5 5781.171296796797u,1.5 5781.172296796797u,0 5782.148836836836u,0 5782.149836836837u,1.5 5783.126376876877u,1.5 5783.127376876877u,0 5788.991617117117u,0 5788.992617117117u,1.5 5789.9691571571575u,1.5 5789.970157157158u,0 5790.946697197197u,0 5790.947697197197u,1.5 5792.901777277278u,1.5 5792.902777277278u,0 5793.879317317317u,0 5793.880317317317u,1.5 5800.722097597598u,1.5 5800.723097597598u,0 5801.699637637637u,0 5801.700637637638u,1.5 5802.677177677678u,1.5 5802.678177677678u,0 5813.430118118118u,0 5813.431118118118u,1.5 5815.385198198198u,1.5 5815.386198198198u,0 5816.362738238237u,0 5816.363738238238u,1.5 5825.160598598599u,1.5 5825.161598598599u,0 5827.115678678679u,0 5827.116678678679u,1.5 5829.070758758759u,1.5 5829.07175875876u,0 5837.868619119119u,0 5837.869619119119u,1.5 5838.8461591591595u,1.5 5838.84715915916u,0 5840.801239239238u,0 5840.802239239239u,1.5 5849.5990995996u,1.5 5849.6000995996u,0 5851.55417967968u,0 5851.55517967968u,1.5 5852.531719719719u,1.5 5852.532719719719u,0 5859.3745u,0 5859.3755u,1.5 5860.352040040039u,1.5 5860.35304004004u,0 5862.30712012012u,0 5862.30812012012u,1.5 5863.2846601601605u,1.5 5863.285660160161u,0 5864.2622002002u,0 5864.2632002002u,1.5 5876.97022072072u,1.5 5876.97122072072u,0 5877.947760760761u,0 5877.948760760762u,1.5 5878.925300800801u,1.5 5878.926300800801u,0 5880.880380880881u,0 5880.881380880881u,1.5 5882.835460960961u,1.5 5882.836460960962u,0 5888.700701201201u,0 5888.701701201201u,1.5 5889.67824124124u,1.5 5889.679241241241u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5899.453641641641u,1.5 5899.4546416416415u,0 5900.431181681682u,0 5900.432181681682u,1.5 5908.251502002002u,1.5 5908.252502002002u,0 5909.229042042041u,0 5909.2300420420415u,1.5 5910.206582082082u,1.5 5910.207582082082u,0 5911.184122122122u,0 5911.185122122122u,1.5 5912.161662162162u,1.5 5912.162662162163u,0 5932.690003003003u,0 5932.691003003003u,1.5 5933.667543043042u,1.5 5933.6685430430425u,0 5935.622623123123u,0 5935.623623123123u,1.5 5936.600163163163u,1.5 5936.601163163164u,0 5938.555243243242u,0 5938.5562432432425u,1.5 5958.106044044043u,1.5 5958.1070440440435u,0 5959.083584084084u,0 5959.084584084084u,1.5 5960.061124124124u,1.5 5960.062124124124u,0 5961.038664164164u,0 5961.039664164165u,1.5 5963.971284284285u,1.5 5963.972284284285u,0 5964.948824324324u,0 5964.949824324324u,1.5 5968.858984484485u,1.5 5968.859984484485u,0 5970.814064564564u,0 5970.815064564565u,1.5 5971.791604604605u,1.5 5971.792604604605u,0 5972.769144644644u,0 5972.7701446446445u,1.5 5973.746684684685u,1.5 5973.747684684685u,0 5979.611924924925u,0 5979.612924924925u,1.5 5980.589464964965u,1.5 5980.590464964966u,0 5983.522085085086u,0 5983.523085085086u,1.5 5984.499625125125u,1.5 5984.500625125125u,0 6006.005506006006u,0 6006.006506006006u,1.5 6006.983046046045u,1.5 6006.9840460460455u,0 6012.848286286287u,0 6012.849286286287u,1.5 6013.825826326326u,1.5 6013.826826326326u,0 6017.735986486487u,0 6017.736986486487u,1.5 6018.713526526526u,1.5 6018.714526526526u,0 6023.601226726726u,0 6023.602226726726u,1.5 6024.578766766767u,1.5 6024.5797667667675u,0 6028.488926926927u,0 6028.489926926927u,1.5 6029.466466966967u,1.5 6029.467466966968u,0 6030.444007007007u,0 6030.445007007007u,1.5 6032.3990870870875u,1.5 6032.400087087088u,0 6033.376627127127u,0 6033.377627127127u,1.5 6036.309247247247u,1.5 6036.310247247247u,0 6037.286787287288u,0 6037.287787287288u,1.5 6055.860048048047u,1.5 6055.861048048047u,0 6056.8375880880885u,0 6056.838588088089u,1.5 6059.770208208208u,1.5 6059.771208208208u,0 6060.747748248248u,0 6060.748748248248u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6068.568068568568u,0 6068.569068568569u,1.5 6070.523148648648u,1.5 6070.524148648648u,0 6071.500688688689u,0 6071.501688688689u,1.5 6072.478228728728u,1.5 6072.479228728728u,0 6074.433308808809u,0 6074.434308808809u,1.5 6075.410848848848u,1.5 6075.411848848848u,0 6087.141329329329u,0 6087.142329329329u,1.5 6088.118869369369u,1.5 6088.11986936937u,0 6090.073949449449u,0 6090.074949449449u,1.5 6101.80442992993u,1.5 6101.80542992993u,0 6102.78196996997u,0 6102.7829699699705u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6106.69213013013u,1.5 6106.69313013013u,0 6107.66967017017u,0 6107.6706701701705u,1.5 6108.64721021021u,1.5 6108.64821021021u,0 6118.422610610611u,0 6118.423610610611u,1.5 6119.40015065065u,1.5 6119.40115065065u,0 6120.3776906906905u,0 6120.378690690691u,1.5 6136.018331331331u,1.5 6136.019331331331u,0 6137.973411411411u,0 6137.974411411411u,1.5 6138.950951451451u,1.5 6138.951951451451u,0 6139.9284914914915u,0 6139.929491491492u,1.5 6140.906031531531u,1.5 6140.907031531531u,0 6147.748811811812u,0 6147.749811811812u,1.5 6148.726351851851u,1.5 6148.727351851851u,0 6151.658971971972u,0 6151.6599719719725u,1.5 6152.636512012012u,1.5 6152.637512012012u,0 6153.614052052051u,0 6153.615052052051u,1.5 6159.4792922922925u,1.5 6159.480292292293u,0 6160.456832332332u,0 6160.457832332332u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6172.187312812813u,0 6172.188312812813u,1.5 6173.164852852852u,1.5 6173.165852852852u,0 6175.119932932933u,0 6175.120932932933u,1.5 6176.097472972973u,1.5 6176.0984729729735u,0 6177.075013013013u,0 6177.076013013013u,1.5 6184.895333333333u,1.5 6184.896333333333u,0 6185.872873373373u,0 6185.8738733733735u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6197.603353853853u,0 6197.604353853853u,1.5 6200.535973973974u,1.5 6200.536973973974u,0 6201.513514014014u,0 6201.514514014014u,1.5 6208.3562942942945u,1.5 6208.357294294295u,0 6215.199074574574u,0 6215.2000745745745u,1.5 6216.176614614615u,1.5 6216.177614614615u,0 6219.109234734734u,0 6219.110234734734u,1.5 6220.086774774775u,1.5 6220.087774774775u,0 6221.064314814815u,0 6221.065314814815u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6231.817255255255u,0 6231.818255255255u,1.5 6232.794795295295u,1.5 6232.795795295296u,0 6239.637575575575u,0 6239.6385755755755u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6256.255756256256u,0 6256.256756256256u,1.5 6257.233296296296u,1.5 6257.234296296297u,0 6260.165916416417u,0 6260.166916416417u,1.5 6261.143456456457u,1.5 6261.144456456457u,0 6262.120996496496u,0 6262.121996496497u,1.5 6268.963776776777u,1.5 6268.964776776777u,0 6269.941316816817u,0 6269.942316816817u,1.5 6270.918856856857u,1.5 6270.919856856857u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6272.873936936937u,1.5 6272.874936936937u,0 6278.739177177177u,0 6278.740177177177u,1.5 6279.716717217217u,1.5 6279.717717217217u,0 6282.649337337337u,0 6282.650337337337u,1.5 6283.626877377377u,1.5 6283.627877377377u,0 6284.604417417418u,0 6284.605417417418u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6291.447197697697u,1.5 6291.448197697698u,0 6304.155218218218u,0 6304.156218218218u,1.5 6305.132758258259u,1.5 6305.133758258259u,0 6306.110298298298u,0 6306.111298298299u,1.5 6307.087838338338u,1.5 6307.088838338338u,0 6308.065378378378u,0 6308.066378378378u,1.5 6313.930618618619u,1.5 6313.931618618619u,0 6314.908158658659u,0 6314.909158658659u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6317.840778778779u,0 6317.841778778779u,1.5 6318.818318818819u,1.5 6318.819318818819u,0 6326.638639139139u,0 6326.639639139139u,1.5 6337.391579579579u,1.5 6337.392579579579u,0 6339.34665965966u,0 6339.34765965966u,1.5 6340.324199699699u,1.5 6340.3251996997u,0 6342.27927977978u,0 6342.28027977978u,1.5 6343.25681981982u,1.5 6343.25781981982u,0 6350.0996001001u,0 6350.100600100101u,1.5 6351.07714014014u,1.5 6351.07814014014u,0 6352.05468018018u,0 6352.05568018018u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6363.785160660661u,1.5 6363.786160660661u,0 6379.425801301301u,0 6379.426801301302u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6406.7969224224225u,0 6406.797922422423u,1.5 6407.774462462463u,1.5 6407.775462462463u,0 6410.707082582582u,0 6410.708082582582u,1.5 6411.684622622623u,1.5 6411.685622622623u,0 6414.617242742742u,0 6414.618242742742u,1.5 6416.572322822823u,1.5 6416.573322822823u,0 6417.549862862863u,0 6417.550862862863u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6437.100663663664u,1.5 6437.101663663664u,0 6446.876064064064u,0 6446.877064064064u,1.5 6447.853604104104u,1.5 6447.8546041041045u,0 6463.494244744744u,0 6463.495244744744u,1.5 6464.471784784785u,1.5 6464.472784784785u,0 6465.4493248248245u,0 6465.450324824825u,1.5 6466.426864864865u,1.5 6466.427864864865u,0 6468.381944944945u,0 6468.382944944945u,1.5 6469.359484984985u,1.5 6469.360484984985u,0 6471.314565065065u,0 6471.315565065065u,1.5 6472.292105105105u,1.5 6472.2931051051055u,0 6474.247185185185u,0 6474.248185185185u,1.5 6476.202265265266u,1.5 6476.203265265266u,0 6477.179805305305u,0 6477.1808053053055u,1.5 6484.022585585586u,1.5 6484.023585585586u,0 6485.0001256256255u,0 6485.001125625626u,1.5 6488.910285785786u,1.5 6488.911285785786u,0 6489.8878258258255u,0 6489.888825825826u,1.5 6500.640766266267u,1.5 6500.641766266267u,0 6501.618306306306u,0 6501.6193063063065u,1.5 6511.393706706706u,1.5 6511.3947067067065u,0 6512.371246746747u,0 6512.372246746747u,1.5 6517.258946946947u,1.5 6517.259946946947u,0 6518.236486986987u,0 6518.237486986987u,1.5 6520.191567067067u,1.5 6520.192567067067u,0 6521.169107107107u,0 6521.1701071071075u,1.5 6525.079267267268u,1.5 6525.080267267268u,0 6527.034347347347u,0 6527.035347347347u,1.5 6528.9894274274275u,1.5 6528.990427427428u,0 6532.899587587588u,0 6532.900587587588u,1.5 6533.8771276276275u,1.5 6533.878127627628u,0 6535.832207707707u,0 6535.8332077077075u,1.5 6536.809747747748u,1.5 6536.810747747748u,0 6562.225788788789u,0 6562.226788788789u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6565.158408908908u,1.5 6565.1594089089085u,0 6566.135948948949u,0 6566.136948948949u,1.5 6568.0910290290285u,1.5 6568.092029029029u,0 6569.068569069069u,0 6569.069569069069u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.001189189189u,0 6572.002189189189u,1.5 6586.66428978979u,1.5 6586.66528978979u,0 6587.6418298298295u,0 6587.64282982983u,1.5 6588.61936986987u,1.5 6588.62036986987u,0 6590.57444994995u,0 6590.57544994995u,1.5 6591.55198998999u,1.5 6591.55298998999u,0 6600.34985035035u,0 6600.35085035035u,1.5 6601.32739039039u,1.5 6601.32839039039u,0 6604.26001051051u,0 6604.2610105105105u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6607.19263063063u,0 6607.193630630631u,1.5 6618.923111111111u,1.5 6618.924111111111u,0 6619.900651151151u,0 6619.901651151151u,1.5 6621.8557312312305u,1.5 6621.856731231231u,0 6623.810811311311u,0 6623.811811311311u,1.5 6624.788351351351u,1.5 6624.789351351351u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6637.496371871872u,0 6637.497371871872u,1.5 6638.473911911911u,1.5 6638.4749119119115u,0 6639.451451951952u,0 6639.452451951952u,1.5 6649.226852352352u,1.5 6649.227852352352u,0 6650.204392392392u,0 6650.205392392392u,1.5 6651.181932432432u,1.5 6651.182932432433u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6664.867492992993u,1.5 6664.868492992993u,0 6665.845033033032u,0 6665.846033033033u,1.5 6672.687813313313u,1.5 6672.688813313313u,0 6673.665353353353u,0 6673.666353353353u,1.5 6674.642893393393u,1.5 6674.643893393393u,0 6676.597973473474u,0 6676.598973473474u,1.5 6677.575513513513u,1.5 6677.576513513513u,0 6685.395833833833u,0 6685.396833833834u,1.5 6693.216154154154u,1.5 6693.217154154154u,0 6694.193694194194u,0 6694.194694194194u,1.5 6698.103854354354u,1.5 6698.104854354354u,0 6705.924174674675u,0 6705.925174674675u,1.5 6706.901714714714u,1.5 6706.902714714714u,0 6707.879254754755u,0 6707.880254754755u,1.5 6708.856794794795u,1.5 6708.857794794795u,0 6709.834334834834u,0 6709.835334834835u,1.5 6718.632195195195u,1.5 6718.633195195195u,0 6719.609735235234u,0 6719.610735235235u,1.5 6720.587275275276u,1.5 6720.588275275276u,0 6726.452515515515u,0 6726.453515515515u,1.5 6727.430055555555u,1.5 6727.431055555555u,0 6729.385135635635u,0 6729.386135635636u,1.5 6741.115616116116u,1.5 6741.116616116116u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6752.846096596597u,0 6752.847096596597u,1.5 6761.6439569569575u,1.5 6761.644956956958u,0 6768.486737237236u,0 6768.487737237237u,1.5 6769.464277277278u,1.5 6769.465277277278u,0 6771.4193573573575u,0 6771.420357357358u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6780.217217717717u,1.5 6780.218217717717u,0 6782.172297797798u,0 6782.173297797798u,1.5 6783.149837837837u,1.5 6783.150837837838u,0 6791.947698198198u,0 6791.948698198198u,1.5 6802.700638638638u,1.5 6802.7016386386385u,0 6803.678178678679u,0 6803.679178678679u,1.5 6804.655718718718u,1.5 6804.656718718718u,0 6813.453579079079u,0 6813.454579079079u,1.5 6814.431119119119u,1.5 6814.432119119119u,0 6815.4086591591595u,0 6815.40965915916u,1.5 6823.22897947948u,1.5 6823.22997947948u,0 6824.206519519519u,0 6824.207519519519u,1.5 6826.1615995996u,1.5 6826.1625995996u,0 6827.139139639639u,0 6827.1401396396395u,1.5 6828.11667967968u,1.5 6828.11767967968u,0 6835.937u,0 6835.938u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6839.8471601601605u,0 6839.848160160161u,1.5 6848.64502052052u,1.5 6848.64602052052u,0 6849.6225605605605u,0 6849.623560560561u,1.5 6851.57764064064u,1.5 6851.5786406406405u,0 6854.510260760761u,0 6854.511260760762u,1.5 6855.487800800801u,1.5 6855.488800800801u,0 6860.375501001001u,0 6860.376501001001u,1.5 6861.35304104104u,1.5 6861.354041041041u,0 6864.285661161161u,0 6864.286661161162u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6867.218281281282u,0 6867.219281281282u,1.5 6876.016141641641u,1.5 6876.0171416416415u,0 6876.993681681682u,0 6876.994681681682u,1.5 6878.948761761762u,1.5 6878.949761761763u,0 6892.634322322322u,0 6892.635322322322u,1.5 6893.611862362362u,1.5 6893.612862362363u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5 6908.274962962963u,1.5 6908.275962962964u,0 6909.252503003003u,0 6909.253503003003u,1.5 6912.185123123123u,1.5 6912.186123123123u,0 6913.162663163163u,0 6913.163663163164u,1.5 6914.140203203203u,1.5 6914.141203203203u,0 6932.713463963964u,0 6932.714463963965u,1.5 6933.691004004004u,1.5 6933.692004004004u,0 6934.668544044043u,0 6934.6695440440435u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6936.623624124124u,0 6936.624624124124u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6939.556244244243u,0 6939.5572442442435u,1.5 6942.488864364364u,1.5 6942.489864364365u,0 6943.466404404404u,0 6943.467404404404u,1.5 6962.039665165165u,1.5 6962.040665165166u,0 6963.017205205205u,0 6963.018205205205u,1.5 6963.994745245244u,1.5 6963.9957452452445u,0 6964.972285285286u,0 6964.973285285286u,1.5 6967.904905405405u,1.5 6967.905905405405u,0 6968.882445445445u,0 6968.883445445445u,1.5 6969.859985485486u,1.5 6969.860985485486u,0 6970.837525525525u,0 6970.838525525525u,1.5 6971.815065565565u,1.5 6971.816065565566u,0 6972.792605605606u,0 6972.793605605606u,1.5 6973.770145645645u,1.5 6973.771145645645u,0 6974.747685685686u,0 6974.748685685686u,1.5 6976.702765765766u,1.5 6976.703765765767u,0 6978.657845845845u,0 6978.6588458458455u,1.5 6979.635385885886u,1.5 6979.636385885886u,0 6981.590465965966u,0 6981.591465965967u,1.5 6982.568006006006u,1.5 6982.569006006006u,0 6986.478166166166u,0 6986.479166166167u,1.5 6987.455706206206u,1.5 6987.456706206206u,0 6989.410786286287u,0 6989.411786286287u,1.5 6990.388326326326u,1.5 6990.389326326326u,0 6991.365866366366u,0 6991.366866366367u,1.5 6992.343406406406u,1.5 6992.344406406406u,0 6994.298486486487u,0 6994.299486486487u,1.5 6995.276026526526u,1.5 6995.277026526526u,0
vb13 b13 0 pwl 0,0  58.6519024024024u,0 58.652902402402404u,1.5 59.62944244244244u,1.5 59.630442442442444u,0 63.539602602602606u,0 63.54060260260261u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 104.59628428428428u,1.5 104.59728428428429u,0 106.55136436436436u,0 106.55236436436437u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 109.48398448448448u,0 109.48498448448449u,1.5 110.46152452452452u,1.5 110.46252452452453u,0 135.8775655655656u,0 135.87856556556557u,1.5 136.85510560560562u,1.5 136.8561056056056u,0 137.83264564564567u,0 137.83364564564565u,1.5 158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 164.22622672672674u,1.5 164.2272267267267u,0 184.7545675675676u,0 184.75556756756757u,1.5 185.73210760760762u,1.5 185.7331076076076u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 188.66472772772775u,0 188.66572772772773u,1.5 207.2379884884885u,1.5 207.23898848848847u,0 208.21552852852852u,0 208.2165285285285u,1.5 210.17060860860863u,1.5 210.1716086086086u,0 229.72140940940943u,0 229.7224094094094u,1.5 230.69894944944946u,1.5 230.69994944944943u,0 231.6764894894895u,0 231.6774894894895u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 270.77809109109114u,0 270.7790910910911u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 272.73317117117114u,0 272.7341711711711u,1.5 289.35135185185186u,1.5 289.35235185185184u,0 290.32889189189194u,0 290.3298918918919u,1.5 294.23905205205205u,1.5 294.240052052052u,0 313.78985285285285u,0 313.7908528528528u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 315.74493293293295u,0 315.74593293293293u,1.5 317.700013013013u,1.5 317.701013013013u,0 318.67755305305303u,0 318.678553053053u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 336.2732737737738u,0 336.27427377377376u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 338.2283538538539u,0 338.22935385385387u,1.5 340.18343393393394u,1.5 340.1844339339339u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 389.06043593593597u,1.5 389.06143593593595u,0 390.037975975976u,0 390.038975975976u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 395.90321621621626u,1.5 395.90421621621624u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 432.07219769769773u,0 432.0731976976977u,1.5 433.04973773773776u,1.5 433.05073773773773u,0 434.0272777777778u,0 434.02827777777776u,1.5 435.00481781781787u,1.5 435.00581781781784u,0 435.98235785785783u,0 435.9833578578578u,1.5 437.93743793793794u,1.5 437.9384379379379u,0 438.91497797797797u,0 438.91597797797795u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 561.107482982983u,0 561.108482982983u,1.5 563.0625630630631u,1.5 563.063563063063u,0 564.0401031031031u,0 564.0411031031031u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 568.9278033033033u,0 568.9288033033033u,1.5 569.9053433433434u,1.5 569.9063433433433u,0 602.1641646646647u,0 602.1651646646646u,1.5 603.1417047047047u,1.5 603.1427047047047u,0 605.0967847847849u,0 605.0977847847848u,1.5 606.0743248248249u,1.5 606.0753248248249u,0 607.0518648648649u,0 607.0528648648649u,1.5 637.355606106106u,1.5 637.356606106106u,0 660.816567067067u,0 660.817567067067u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 662.7716471471472u,0 662.7726471471472u,1.5 663.7491871871872u,1.5 663.7501871871872u,0 664.7267272272272u,0 664.7277272272272u,1.5 685.255068068068u,1.5 685.256068068068u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 707.7384889889889u,0 707.7394889889889u,1.5 708.716029029029u,1.5 708.7170290290289u,0 709.693569069069u,0 709.694569069069u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 729.24436986987u,1.5 729.2453698698699u,0 730.22190990991u,0 730.22290990991u,1.5 731.19944994995u,1.5 731.20044994995u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 771.2785915915915u,0 771.2795915915915u,1.5 772.2561316316315u,1.5 772.2571316316315u,0 790.8293923923924u,0 790.8303923923924u,1.5 792.7844724724725u,1.5 792.7854724724725u,0 793.7620125125126u,0 793.7630125125125u,1.5 814.2903533533533u,1.5 814.2913533533533u,0 815.2678933933934u,0 815.2688933933933u,1.5 816.2454334334335u,1.5 816.2464334334335u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 841.6614744744745u,0 841.6624744744745u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 868.0550555555556u,0 868.0560555555555u,1.5 869.0325955955957u,1.5 869.0335955955957u,0 894.4486366366367u,0 894.4496366366367u,1.5 896.4037167167166u,1.5 896.4047167167166u,0 897.3812567567567u,0 897.3822567567566u,1.5 927.684997997998u,1.5 927.685997997998u,0 928.6625380380381u,0 928.663538038038u,1.5 932.5726981981983u,1.5 932.5736981981983u,0 933.5502382382382u,0 933.5512382382382u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 938.4379384384384u,0 938.4389384384384u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 1057.6978233233233u,0 1057.6988233233235u,1.5 1058.6753633633632u,1.5 1058.6763633633634u,0 1061.6079834834834u,0 1061.6089834834836u,1.5 1062.5855235235235u,1.5 1062.5865235235237u,0 1065.5181436436435u,0 1065.5191436436437u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1070.4058438438437u,1.5 1070.406843843844u,0 1071.3833838838837u,0 1071.3843838838839u,1.5 1102.6646651651652u,1.5 1102.6656651651654u,0 1103.642205205205u,0 1103.6432052052053u,1.5 1104.6197452452452u,1.5 1104.6207452452454u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1107.5523653653654u,1.5 1107.5533653653656u,0 1108.5299054054053u,0 1108.5309054054055u,1.5 1109.5074454454455u,1.5 1109.5084454454457u,0 1134.9234864864864u,0 1134.9244864864866u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1161.3170675675676u,1.5 1161.3180675675678u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1163.2721476476477u,1.5 1163.2731476476479u,0 1164.2496876876876u,0 1164.2506876876878u,1.5 1165.2272277277275u,1.5 1165.2282277277277u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1208.2389894894895u,0 1208.2399894894897u,1.5 1210.1940695695696u,1.5 1210.1950695695698u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1231.6999504504504u,0 1231.7009504504506u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1254.1833713713713u,1.5 1254.1843713713715u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1269.8240120120117u,1.5 1269.825012012012u,0 1270.8015520520519u,0 1270.802552052052u,1.5 1271.779092092092u,1.5 1271.7800920920922u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1291.3298928928928u,0 1291.330892892893u,1.5 1292.3074329329327u,1.5 1292.3084329329329u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1315.7683938938937u,1.5 1315.769393893894u,0 1316.7459339339337u,0 1316.7469339339339u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1342.1619749749748u,1.5 1342.162974974975u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1367.578016016016u,1.5 1367.579016016016u,0 1368.5555560560558u,0 1368.556556056056u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1400.8143773773772u,0 1400.8153773773774u,1.5 1401.7919174174174u,1.5 1401.7929174174176u,0 1431.1181186186186u,0 1431.1191186186188u,1.5 1432.0956586586585u,1.5 1432.0966586586587u,0 1433.0731986986987u,0 1433.0741986986989u,1.5 1434.0507387387386u,1.5 1434.0517387387388u,0 1436.0058188188189u,0 1436.006818818819u,1.5 1438.938438938939u,1.5 1438.9394389389392u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1562.108483983984u,1.5 1562.109483983984u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1565.041104104104u,1.5 1565.0421041041043u,0 1566.996184184184u,0 1566.997184184184u,1.5 1567.973724224224u,1.5 1567.9747242242242u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1603.1651656656657u,1.5 1603.1661656656659u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1607.0753258258258u,0 1607.076325825826u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1662.795108108108u,0 1662.7961081081082u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1689.1886891891893u,0 1689.1896891891895u,1.5 1690.1662292292292u,1.5 1690.1672292292294u,0 1704.8293298298297u,0 1704.83032982983u,1.5 1705.8068698698698u,1.5 1705.80786986987u,0 1707.76194994995u,0 1707.76294994995u,1.5 1728.2902907907908u,1.5 1728.291290790791u,0 1729.2678308308307u,0 1729.268830830831u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1752.7287917917918u,0 1752.729791791792u,1.5 1767.3918923923923u,1.5 1767.3928923923925u,0 1768.3694324324322u,0 1768.3704324324324u,1.5 1771.3020525525524u,1.5 1771.3030525525526u,0 1790.852853353353u,0 1790.8538533533533u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1794.7630135135132u,1.5 1794.7640135135134u,0 1795.7405535535534u,0 1795.7415535535536u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1839.7298553553553u,0 1839.7308553553555u,1.5 1863.1908163163164u,1.5 1863.1918163163166u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1866.1234364364361u,1.5 1866.1244364364363u,0 1889.5843973973974u,0 1889.5853973973976u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1896.4271776776775u,0 1896.4281776776777u,1.5 1897.4047177177176u,1.5 1897.4057177177178u,0 1898.3822577577575u,0 1898.3832577577577u,1.5 1899.3597977977977u,1.5 1899.3607977977979u,0 1900.3373378378376u,0 1900.3383378378378u,1.5 1929.6635390390388u,1.5 1929.664539039039u,0 1930.641079079079u,0 1930.6420790790792u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1940.4164794794794u,0 1940.4174794794797u,1.5 1941.3940195195194u,1.5 1941.3950195195196u,0 1943.3490995995994u,0 1943.3500995995996u,1.5 1944.3266396396396u,1.5 1944.3276396396398u,0 2059.676364364364u,0 2059.677364364364u,1.5 2060.6539044044043u,1.5 2060.6549044044045u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2067.4966846846846u,0 2067.497684684685u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2070.429304804805u,0 2070.430304804805u,1.5 2103.665666166166u,1.5 2103.666666166166u,0 2104.643206206206u,0 2104.644206206206u,1.5 2105.620746246246u,1.5 2105.6217462462464u,0 2134.946947447447u,0 2134.9479474474474u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2137.8795675675674u,0 2137.8805675675676u,1.5 2138.8571076076073u,1.5 2138.8581076076075u,0 2139.8346476476477u,0 2139.835647647648u,1.5 2162.3180685685684u,1.5 2162.3190685685686u,0 2163.2956086086083u,0 2163.2966086086085u,1.5 2164.2731486486487u,1.5 2164.274148648649u,0 2184.8014894894895u,0 2184.8024894894897u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2187.7341096096093u,0 2187.7351096096095u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2227.813251251251u,0 2227.8142512512513u,1.5 2228.790791291291u,1.5 2228.7917912912912u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2230.745871371371u,1.5 2230.746871371371u,0 2231.7234114114112u,0 2231.7244114114114u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2254.2068323323324u,1.5 2254.2078323323326u,0 2268.869932932933u,0 2268.870932932933u,1.5 2269.847472972973u,1.5 2269.848472972973u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2290.3758138138137u,1.5 2290.376813813814u,0 2292.330893893894u,0 2292.331893893894u,1.5 2293.308433933934u,1.5 2293.309433933934u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2314.8143148148147u,1.5 2314.815314814815u,0 2316.769394894895u,0 2316.770394894895u,1.5 2317.746934934935u,1.5 2317.747934934935u,0 2318.724474974975u,0 2318.725474974975u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2340.2303558558556u,0 2340.231355855856u,1.5 2341.207895895896u,1.5 2341.208895895896u,0 2359.7811566566565u,0 2359.7821566566568u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2365.646396896897u,0 2365.647396896897u,1.5 2367.6014769769768u,1.5 2367.602476976977u,0 2368.5790170170167u,0 2368.580017017017u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2397.905218218218u,1.5 2397.9062182182183u,0 2432.119119619619u,0 2432.1201196196193u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2435.05173973974u,1.5 2435.05273973974u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.9843598598595u,1.5 2437.9853598598597u,0 2438.9618998999u,0 2438.9628998999u,1.5 2554.3116246246245u,1.5 2554.3126246246247u,0 2555.2891646646644u,0 2555.2901646646646u,1.5 2558.2217847847846u,1.5 2558.222784784785u,0 2559.1993248248245u,0 2559.2003248248247u,1.5 2560.1768648648645u,1.5 2560.1778648648647u,0 2562.1319449449447u,0 2562.132944944945u,1.5 2565.064565065065u,1.5 2565.065565065065u,0 2566.042105105105u,0 2566.043105105105u,1.5 2567.019645145145u,1.5 2567.0206451451454u,0 2567.997185185185u,0 2567.9981851851853u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2608.0763268268265u,0 2608.0773268268267u,1.5 2634.469907907908u,1.5 2634.470907907908u,0 2635.4474479479477u,0 2635.448447947948u,1.5 2637.402528028028u,1.5 2637.403528028028u,0 2657.9308688688684u,0 2657.9318688688686u,1.5 2658.9084089089088u,1.5 2658.909408908909u,0 2659.8859489489487u,0 2659.886948948949u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2665.751189189189u,1.5 2665.7521891891893u,0 2666.7287292292294u,0 2666.7297292292296u,1.5 2685.30198998999u,1.5 2685.3029899899902u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2689.21215015015u,0 2689.2131501501503u,1.5 2690.18969019019u,1.5 2690.1906901901903u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2710.718031031031u,1.5 2710.719031031031u,0 2711.695571071071u,0 2711.696571071071u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2730.268831831832u,1.5 2730.269831831832u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2750.7971726726723u,0 2750.7981726726725u,1.5 2751.7747127127127u,1.5 2751.775712712713u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2773.2805935935935u,1.5 2773.2815935935937u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2839.753316316316u,1.5 2839.7543163163164u,0 2840.730856356356u,0 2840.7318563563563u,1.5 2860.281657157157u,1.5 2860.2826571571572u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2865.169357357357u,0 2865.1703573573573u,1.5 2866.1468973973974u,1.5 2866.1478973973976u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2930.66454004004u,1.5 2930.66554004004u,0 2931.64208008008u,0 2931.6430800800804u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2938.48486036036u,0 2938.48586036036u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2941.4174804804807u,1.5 2941.418480480481u,0 2942.39502052052u,0 2942.3960205205203u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 3062.6324454454452u,0 3062.6334454454454u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3066.5426056056053u,1.5 3066.5436056056055u,0 3067.5201456456457u,0 3067.521145645646u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3104.666667167167u,0 3104.667667167167u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3135.947948448448u,0 3135.9489484484484u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3207.308371371371u,1.5 3207.309371371371u,0 3227.836712212212u,0 3227.8377122122124u,1.5 3228.814252252252u,1.5 3228.8152522522523u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3232.724412412412u,1.5 3232.7254124124124u,0 3233.701952452452u,0 3233.7029524524523u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3273.781094094094u,0 3273.782094094094u,1.5 3290.3992747747743u,1.5 3290.4002747747745u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3294.309434934935u,1.5 3294.310434934935u,0 3309.9500755755753u,0 3309.9510755755755u,1.5 3310.927615615615u,1.5 3310.9286156156154u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3335.366116616616u,1.5 3335.3671166166164u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3365.6698578578576u,1.5 3365.6708578578578u,0 3366.647397897898u,0 3366.648397897898u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3390.1083588588585u,0 3390.1093588588587u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.996059059059u,0 3394.997059059059u,1.5 3396.9511391391393u,1.5 3396.9521391391395u,0 3431.1650405405403u,0 3431.1660405405405u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3434.0976606606605u,0 3434.0986606606607u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3436.052740740741u,0 3436.053740740741u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.020646146146u,0 3568.0216461461464u,1.5 3568.998186186186u,1.5 3568.9991861861863u,0 3603.2120875875876u,0 3603.213087587588u,1.5 3605.1671676676674u,1.5 3605.1681676676676u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3607.1222477477477u,1.5 3607.123247747748u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3635.4709089089088u,1.5 3635.471908908909u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3637.425988988989u,1.5 3637.4269889889893u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3688.258071071071u,1.5 3688.259071071071u,0 3706.831331831832u,0 3706.832331831832u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3732.2473728728723u,0 3732.2483728728726u,1.5 3733.2249129129127u,1.5 3733.225912912913u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3772.326514514514u,1.5 3772.3275145145144u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3812.405656156156u,1.5 3812.4066561561563u,0 3813.383196196196u,0 3813.384196196196u,1.5 3814.3607362362363u,1.5 3814.3617362362365u,0 3815.338276276276u,0 3815.339276276276u,1.5 3816.315816316316u,1.5 3816.3168163163164u,0 3817.293356356356u,0 3817.2943563563563u,1.5 3818.2708963963964u,1.5 3818.2718963963966u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3836.844157157157u,1.5 3836.8451571571572u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3887.6762392392393u,0 3887.6772392392395u,1.5 3888.653779279279u,1.5 3888.6547792792794u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3895.4965595595595u,0 3895.4975595595597u,1.5 3933.6206211211206u,1.5 3933.621621121121u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3938.508321321321u,0 3938.5093213213213u,1.5 3939.4858613613615u,1.5 3939.4868613613617u,0 4057.768206206206u,0 4057.769206206206u,1.5 4058.7457462462457u,1.5 4058.746746246246u,0 4061.6783663663664u,0 4061.6793663663666u,1.5 4062.6559064064063u,1.5 4062.6569064064065u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4065.588526526526u,1.5 4065.5895265265262u,0 4066.566066566567u,0 4066.567066566567u,1.5 4067.5436066066063u,1.5 4067.5446066066065u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4101.757508008008u,1.5 4101.758508008008u,0 4102.735048048047u,0 4102.736048048047u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4105.667668168168u,0 4105.668668168169u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4134.993869369369u,0 4134.99486936937u,1.5 4137.9264894894895u,1.5 4137.92748948949u,0 4138.904029529529u,0 4138.905029529529u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4183.870871371371u,0 4183.8718713713715u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4209.286912412412u,1.5 4209.287912412412u,0 4225.9050930930935u,0 4225.906093093094u,1.5 4226.882633133133u,1.5 4226.883633133133u,0 4229.815253253253u,0 4229.816253253253u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4268.916854854855u,0 4268.917854854855u,1.5 4270.871934934935u,1.5 4270.872934934935u,0 4272.827015015015u,0 4272.828015015015u,1.5 4289.4451956956955u,1.5 4289.446195695696u,0 4290.422735735735u,0 4290.423735735735u,1.5 4292.377815815816u,1.5 4292.378815815816u,0 4293.355355855856u,0 4293.356355855856u,1.5 4294.3328958958955u,1.5 4294.333895895896u,0 4313.8836966966965u,0 4313.884696696697u,1.5 4336.367117617618u,1.5 4336.368117617618u,0 4337.344657657658u,0 4337.345657657658u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4342.232357857858u,1.5 4342.233357857858u,0 4361.783158658659u,0 4361.784158658659u,1.5 4362.760698698698u,1.5 4362.761698698699u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4368.625938938939u,1.5 4368.626938938939u,0 4369.603478978979u,0 4369.604478978979u,1.5 4390.13181981982u,1.5 4390.13281981982u,0 4391.10935985986u,0 4391.11035985986u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.99706006006u,1.5 4395.99806006006u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4438.031281781782u,0 4438.032281781782u,1.5 4440.963901901901u,1.5 4440.964901901902u,0 4441.941441941942u,0 4441.942441941942u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4566.0890270270265u,0 4566.090027027027u,1.5 4567.066567067067u,1.5 4567.067567067067u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4609.100788788789u,1.5 4609.101788788789u,0 4610.0783288288285u,0 4610.079328828829u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4636.471909909909u,0 4636.4729099099095u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4704.899712712712u,0 4704.900712712712u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4731.293293793794u,0 4731.294293793794u,1.5 4732.270833833833u,1.5 4732.271833833834u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4768.439815315315u,1.5 4768.440815315315u,0 4769.4173553553555u,0 4769.418355355356u,1.5 4771.372435435435u,1.5 4771.373435435436u,0 4793.8558563563565u,0 4793.856856356357u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4840.777778278279u,1.5 4840.778778278279u,0 4841.755318318318u,0 4841.756318318318u,1.5 4863.261199199199u,1.5 4863.262199199199u,0 4864.238739239238u,0 4864.239739239239u,1.5 4866.193819319319u,1.5 4866.194819319319u,0 4891.6098603603605u,0 4891.610860360361u,1.5 4892.5874004004u,1.5 4892.5884004004u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4894.542480480481u,1.5 4894.543480480481u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4898.45264064064u,1.5 4898.4536406406405u,0 4899.430180680681u,0 4899.431180680681u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4938.531782282283u,1.5 4938.532782282283u,0 4940.486862362362u,0 4940.487862362363u,1.5 4941.464402402402u,1.5 4941.465402402402u,0 5057.791667167167u,0 5057.792667167168u,1.5 5058.769207207207u,1.5 5058.770207207207u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5064.634447447447u,0 5064.635447447447u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5135.01733033033u,0 5135.01833033033u,1.5 5135.99487037037u,1.5 5135.9958703703705u,0 5136.97241041041u,0 5136.97341041041u,1.5 5160.433371371371u,1.5 5160.4343713713715u,0 5161.410911411411u,0 5161.411911411411u,1.5 5162.388451451451u,1.5 5162.389451451451u,0 5186.826952452452u,0 5186.827952452452u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5232.771334334334u,0 5232.772334334334u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5271.872935935936u,0 5271.873935935936u,1.5 5289.468656656657u,1.5 5289.469656656657u,0 5290.4461966966965u,0 5290.447196696697u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5294.356356856857u,0 5294.357356856857u,1.5 5295.3338968968965u,1.5 5295.334896896897u,0 5312.929617617618u,0 5312.930617617618u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5337.368118618619u,1.5 5337.369118618619u,0 5338.345658658659u,0 5338.346658658659u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5362.78415965966u,0 5362.78515965966u,1.5 5363.761699699699u,1.5 5363.7626996997u,0 5364.739239739739u,0 5364.740239739739u,1.5 5366.69431981982u,1.5 5366.69531981982u,0 5367.67185985986u,0 5367.67285985986u,1.5 5394.065440940941u,1.5 5394.066440940941u,0 5395.042980980981u,0 5395.043980980981u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5396.998061061061u,0 5396.999061061061u,1.5 5397.975601101101u,1.5 5397.976601101102u,0 5398.953141141141u,0 5398.954141141141u,1.5 5399.930681181181u,1.5 5399.931681181181u,0 5430.2344224224225u,0 5430.235422422423u,1.5 5431.211962462463u,1.5 5431.212962462463u,0 5432.189502502502u,0 5432.190502502503u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5438.054742742742u,1.5 5438.055742742742u,0 5439.032282782783u,0 5439.033282782783u,1.5 5440.009822822823u,1.5 5440.010822822823u,0 5440.987362862863u,0 5440.988362862863u,1.5 5444.897523023023u,1.5 5444.898523023023u,0 5445.875063063063u,0 5445.876063063063u,1.5 5558.292167667668u,1.5 5558.293167667668u,0 5559.269707707707u,0 5559.2707077077075u,1.5 5562.2023278278275u,1.5 5562.203327827828u,0 5563.179867867868u,0 5563.180867867868u,1.5 5566.112487987988u,1.5 5566.113487987988u,0 5567.0900280280275u,0 5567.091028028028u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5570.022648148148u,0 5570.023648148148u,1.5 5571.000188188188u,1.5 5571.001188188188u,0 5600.326389389389u,0 5600.327389389389u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5605.21408958959u,0 5605.21508958959u,1.5 5608.146709709709u,1.5 5608.1477097097095u,0 5609.12424974975u,0 5609.12524974975u,1.5 5633.562750750751u,1.5 5633.563750750751u,0 5634.540290790791u,0 5634.541290790791u,1.5 5636.495370870871u,1.5 5636.496370870871u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5638.450450950951u,1.5 5638.451450950951u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5664.8440320320315u,1.5 5664.845032032032u,0 5665.821572072072u,0 5665.822572072072u,1.5 5682.439752752753u,1.5 5682.440752752753u,0 5683.417292792793u,0 5683.418292792793u,1.5 5685.372372872873u,1.5 5685.373372872873u,0 5688.304992992993u,0 5688.305992992993u,1.5 5689.282533033032u,1.5 5689.283533033033u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5727.406594594595u,1.5 5727.407594594595u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5772.373436436436u,1.5 5772.374436436437u,0 5788.991617117117u,0 5788.992617117117u,1.5 5789.9691571571575u,1.5 5789.970157157158u,0 5790.946697197197u,0 5790.947697197197u,1.5 5792.901777277278u,1.5 5792.902777277278u,0 5793.879317317317u,0 5793.880317317317u,1.5 5813.430118118118u,1.5 5813.431118118118u,0 5815.385198198198u,0 5815.386198198198u,1.5 5816.362738238237u,1.5 5816.363738238238u,0 5837.868619119119u,0 5837.869619119119u,1.5 5838.8461591591595u,1.5 5838.84715915916u,0 5840.801239239238u,0 5840.802239239239u,1.5 5859.3745u,1.5 5859.3755u,0 5860.352040040039u,0 5860.35304004004u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5863.2846601601605u,0 5863.285660160161u,1.5 5864.2622002002u,1.5 5864.2632002002u,0 5888.700701201201u,0 5888.701701201201u,1.5 5889.67824124124u,1.5 5889.679241241241u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5899.453641641641u,1.5 5899.4546416416415u,0 5900.431181681682u,0 5900.432181681682u,1.5 5932.690003003003u,1.5 5932.691003003003u,0 5933.667543043042u,0 5933.6685430430425u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5936.600163163163u,0 5936.601163163164u,1.5 5938.555243243242u,1.5 5938.5562432432425u,0 6055.860048048047u,0 6055.861048048047u,1.5 6056.8375880880885u,1.5 6056.838588088089u,0 6059.770208208208u,0 6059.771208208208u,1.5 6060.747748248248u,1.5 6060.748748248248u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6068.568068568568u,1.5 6068.569068568569u,0 6070.523148648648u,0 6070.524148648648u,1.5 6071.500688688689u,1.5 6071.501688688689u,0 6072.478228728728u,0 6072.479228728728u,1.5 6074.433308808809u,1.5 6074.434308808809u,0 6075.410848848848u,0 6075.411848848848u,1.5 6101.80442992993u,1.5 6101.80542992993u,0 6102.78196996997u,0 6102.7829699699705u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6106.69213013013u,1.5 6106.69313013013u,0 6107.66967017017u,0 6107.6706701701705u,1.5 6108.64721021021u,1.5 6108.64821021021u,0 6136.018331331331u,0 6136.019331331331u,1.5 6137.973411411411u,1.5 6137.974411411411u,0 6138.950951451451u,0 6138.951951451451u,1.5 6139.9284914914915u,1.5 6139.929491491492u,0 6140.906031531531u,0 6140.907031531531u,1.5 6159.4792922922925u,1.5 6159.480292292293u,0 6160.456832332332u,0 6160.457832332332u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6184.895333333333u,0 6184.896333333333u,1.5 6185.872873373373u,1.5 6185.8738733733735u,0 6186.850413413413u,0 6186.851413413413u,1.5 6208.3562942942945u,1.5 6208.357294294295u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6232.794795295295u,0 6232.795795295296u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6268.963776776777u,0 6268.964776776777u,1.5 6269.941316816817u,1.5 6269.942316816817u,0 6270.918856856857u,0 6270.919856856857u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6272.873936936937u,0 6272.874936936937u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6291.447197697697u,1.5 6291.448197697698u,0 6313.930618618619u,0 6313.931618618619u,1.5 6314.908158658659u,1.5 6314.909158658659u,0 6315.885698698698u,0 6315.886698698699u,1.5 6317.840778778779u,1.5 6317.841778778779u,0 6318.818318818819u,0 6318.819318818819u,1.5 6337.391579579579u,1.5 6337.392579579579u,0 6339.34665965966u,0 6339.34765965966u,1.5 6340.324199699699u,1.5 6340.3251996997u,0 6342.27927977978u,0 6342.28027977978u,1.5 6343.25681981982u,1.5 6343.25781981982u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6363.785160660661u,0 6363.786160660661u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6437.100663663664u,0 6437.101663663664u,1.5 6446.876064064064u,1.5 6446.877064064064u,0 6447.853604104104u,0 6447.8546041041045u,1.5 6562.225788788789u,1.5 6562.226788788789u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6565.158408908908u,0 6565.1594089089085u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6568.0910290290285u,0 6568.092029029029u,1.5 6569.068569069069u,1.5 6569.069569069069u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.001189189189u,1.5 6572.002189189189u,0 6600.34985035035u,0 6600.35085035035u,1.5 6601.32739039039u,1.5 6601.32839039039u,0 6604.26001051051u,0 6604.2610105105105u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6607.19263063063u,0 6607.193630630631u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6637.496371871872u,1.5 6637.497371871872u,0 6638.473911911911u,0 6638.4749119119115u,1.5 6639.451451951952u,1.5 6639.452451951952u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6664.867492992993u,1.5 6664.868492992993u,0 6665.845033033032u,0 6665.846033033033u,1.5 6685.395833833833u,1.5 6685.396833833834u,0 6705.924174674675u,0 6705.925174674675u,1.5 6706.901714714714u,1.5 6706.902714714714u,0 6707.879254754755u,0 6707.880254754755u,1.5 6708.856794794795u,1.5 6708.857794794795u,0 6709.834334834834u,0 6709.835334834835u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6727.430055555555u,0 6727.431055555555u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6752.846096596597u,0 6752.847096596597u,1.5 6768.486737237236u,1.5 6768.487737237237u,0 6769.464277277278u,0 6769.465277277278u,1.5 6771.4193573573575u,1.5 6771.420357357358u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6791.947698198198u,0 6791.948698198198u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6814.431119119119u,0 6814.432119119119u,1.5 6815.4086591591595u,1.5 6815.40965915916u,0 6835.937u,0 6835.938u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6839.8471601601605u,0 6839.848160160161u,1.5 6860.375501001001u,1.5 6860.376501001001u,0 6861.35304104104u,0 6861.354041041041u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6866.24074124124u,0 6866.241741241241u,1.5 6867.218281281282u,1.5 6867.219281281282u,0 6892.634322322322u,0 6892.635322322322u,1.5 6893.611862362362u,1.5 6893.612862362363u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5 6932.713463963964u,1.5 6932.714463963965u,0 6933.691004004004u,0 6933.692004004004u,1.5 6934.668544044043u,1.5 6934.6695440440435u,0 6935.646084084084u,0 6935.647084084084u,1.5 6936.623624124124u,1.5 6936.624624124124u,0 6938.578704204204u,0 6938.579704204204u,1.5 6939.556244244243u,1.5 6939.5572442442435u,0 6942.488864364364u,0 6942.489864364365u,1.5 6943.466404404404u,1.5 6943.467404404404u,0
vb14 b14 0 pwl 0,0  104.59628428428428u,0 104.59728428428429u,1.5 106.55136436436436u,1.5 106.55236436436437u,0 107.5289044044044u,0 107.5299044044044u,1.5 109.48398448448448u,1.5 109.48498448448449u,0 110.46152452452452u,0 110.46252452452453u,1.5 158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 164.22622672672674u,1.5 164.2272267267267u,0 207.2379884884885u,0 207.23898848848847u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 210.17060860860863u,0 210.1716086086086u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 289.35135185185186u,0 289.35235185185184u,1.5 290.32889189189194u,1.5 290.3298918918919u,0 294.23905205205205u,0 294.240052052052u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 336.2732737737738u,0 336.27427377377376u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 338.2283538538539u,0 338.22935385385387u,1.5 340.18343393393394u,1.5 340.1844339339339u,0 389.06043593593597u,0 389.06143593593595u,1.5 390.037975975976u,1.5 390.038975975976u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 395.90321621621626u,0 395.90421621621624u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 602.1641646646647u,1.5 602.1651646646646u,0 603.1417047047047u,0 603.1427047047047u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 606.0743248248249u,0 606.0753248248249u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 660.816567067067u,0 660.817567067067u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 662.7716471471472u,0 662.7726471471472u,1.5 663.7491871871872u,1.5 663.7501871871872u,0 664.7267272272272u,0 664.7277272272272u,1.5 707.7384889889889u,1.5 707.7394889889889u,0 708.716029029029u,0 708.7170290290289u,1.5 709.693569069069u,1.5 709.694569069069u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 790.8293923923924u,1.5 790.8303923923924u,0 792.7844724724725u,0 792.7854724724725u,1.5 793.7620125125126u,1.5 793.7630125125125u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 841.6614744744745u,0 841.6624744744745u,1.5 894.4486366366367u,1.5 894.4496366366367u,0 896.4037167167166u,0 896.4047167167166u,1.5 897.3812567567567u,1.5 897.3822567567566u,0 1102.6646651651652u,0 1102.6656651651654u,1.5 1103.642205205205u,1.5 1103.6432052052053u,0 1104.6197452452452u,0 1104.6207452452454u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1107.5523653653654u,0 1107.5533653653656u,1.5 1108.5299054054053u,1.5 1108.5309054054055u,0 1109.5074454454455u,0 1109.5084454454457u,1.5 1161.3170675675676u,1.5 1161.3180675675678u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1163.2721476476477u,1.5 1163.2731476476479u,0 1164.2496876876876u,0 1164.2506876876878u,1.5 1165.2272277277275u,1.5 1165.2282277277277u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1208.2389894894895u,1.5 1208.2399894894897u,0 1210.1940695695696u,0 1210.1950695695698u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1254.1833713713713u,1.5 1254.1843713713715u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1291.3298928928928u,1.5 1291.330892892893u,0 1292.3074329329327u,0 1292.3084329329329u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1342.1619749749748u,1.5 1342.162974974975u,0 1392.016517017017u,0 1392.017517017017u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1400.8143773773772u,1.5 1400.8153773773774u,0 1401.7919174174174u,0 1401.7929174174176u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1603.1651656656657u,0 1603.1661656656659u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1607.0753258258258u,1.5 1607.076325825826u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1662.795108108108u,0 1662.7961081081082u,1.5 1704.8293298298297u,1.5 1704.83032982983u,0 1705.8068698698698u,0 1705.80786986987u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1752.7287917917918u,0 1752.729791791792u,1.5 1790.852853353353u,1.5 1790.8538533533533u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1794.7630135135132u,0 1794.7640135135134u,1.5 1795.7405535535534u,1.5 1795.7415535535536u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1839.7298553553553u,0 1839.7308553553555u,1.5 1889.5843973973974u,1.5 1889.5853973973976u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1896.4271776776775u,1.5 1896.4281776776777u,0 1897.4047177177176u,0 1897.4057177177178u,1.5 1898.3822577577575u,1.5 1898.3832577577577u,0 1899.3597977977977u,0 1899.3607977977979u,1.5 1900.3373378378376u,1.5 1900.3383378378378u,0 2103.665666166166u,0 2103.666666166166u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2105.620746246246u,0 2105.6217462462464u,1.5 2162.3180685685684u,1.5 2162.3190685685686u,0 2163.2956086086083u,0 2163.2966086086085u,1.5 2164.2731486486487u,1.5 2164.274148648649u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2254.2068323323324u,1.5 2254.2078323323326u,0 2290.3758138138137u,0 2290.376813813814u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2293.308433933934u,0 2293.309433933934u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2340.2303558558556u,0 2340.231355855856u,1.5 2341.207895895896u,1.5 2341.208895895896u,0 2393.995058058058u,0 2393.996058058058u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2397.905218218218u,0 2397.9062182182183u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2608.0763268268265u,1.5 2608.0773268268267u,0 2657.9308688688684u,0 2657.9318688688686u,1.5 2658.9084089089088u,1.5 2658.909408908909u,0 2659.8859489489487u,0 2659.886948948949u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2665.751189189189u,1.5 2665.7521891891893u,0 2666.7287292292294u,0 2666.7297292292296u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2710.718031031031u,0 2710.719031031031u,1.5 2711.695571071071u,1.5 2711.696571071071u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2750.7971726726723u,0 2750.7981726726725u,1.5 2751.7747127127127u,1.5 2751.775712712713u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2839.753316316316u,1.5 2839.7543163163164u,0 2840.730856356356u,0 2840.7318563563563u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 3103.689127127127u,0 3103.690127127127u,1.5 3104.666667167167u,1.5 3104.667667167167u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3207.308371371371u,0 3207.309371371371u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3290.3992747747743u,0 3290.4002747747745u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3294.309434934935u,0 3294.310434934935u,1.5 3335.366116616616u,1.5 3335.3671166166164u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3390.1083588588585u,1.5 3390.1093588588587u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3396.9511391391393u,0 3396.9521391391395u,1.5 3603.2120875875876u,1.5 3603.213087587588u,0 3605.1671676676674u,0 3605.1681676676676u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3607.1222477477477u,0 3607.123247747748u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3706.831331831832u,1.5 3706.832331831832u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3836.844157157157u,1.5 3836.8451571571572u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 3887.6762392392393u,1.5 3887.6772392392395u,0 3888.653779279279u,0 3888.6547792792794u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3895.4965595595595u,1.5 3895.4975595595597u,0 4101.757508008008u,0 4101.758508008008u,1.5 4102.735048048047u,1.5 4102.736048048047u,0 4104.690128128128u,0 4104.691128128128u,1.5 4105.667668168168u,1.5 4105.668668168169u,0 4106.645208208208u,0 4106.646208208208u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4209.286912412412u,0 4209.287912412412u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4289.4451956956955u,0 4289.446195695696u,1.5 4290.422735735735u,1.5 4290.423735735735u,0 4292.377815815816u,0 4292.378815815816u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4294.3328958958955u,0 4294.333895895896u,1.5 4336.367117617618u,1.5 4336.368117617618u,0 4337.344657657658u,0 4337.345657657658u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4342.232357857858u,1.5 4342.233357857858u,0 4390.13181981982u,0 4390.13281981982u,1.5 4391.10935985986u,1.5 4391.11035985986u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.99706006006u,0 4395.99806006006u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4609.100788788789u,0 4609.101788788789u,1.5 4610.0783288288285u,1.5 4610.079328828829u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4704.899712712712u,1.5 4704.900712712712u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4793.8558563563565u,1.5 4793.856856356357u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4840.777778278279u,1.5 4840.778778278279u,0 4841.755318318318u,0 4841.756318318318u,1.5 4891.6098603603605u,1.5 4891.610860360361u,0 4892.5874004004u,0 4892.5884004004u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4894.542480480481u,0 4894.543480480481u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4898.45264064064u,0 4898.4536406406405u,1.5 4899.430180680681u,1.5 4899.431180680681u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5160.433371371371u,1.5 5160.4343713713715u,0 5161.410911411411u,0 5161.411911411411u,1.5 5162.388451451451u,1.5 5162.389451451451u,0 5208.332833333333u,0 5208.333833333333u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5289.468656656657u,0 5289.469656656657u,1.5 5290.4461966966965u,1.5 5290.447196696697u,0 5292.401276776777u,0 5292.402276776777u,1.5 5294.356356856857u,1.5 5294.357356856857u,0 5295.3338968968965u,0 5295.334896896897u,1.5 5337.368118618619u,1.5 5337.369118618619u,0 5338.345658658659u,0 5338.346658658659u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5394.065440940941u,0 5394.066440940941u,1.5 5395.042980980981u,1.5 5395.043980980981u,0 5396.020521021021u,0 5396.021521021021u,1.5 5396.998061061061u,1.5 5396.999061061061u,0 5397.975601101101u,0 5397.976601101102u,1.5 5398.953141141141u,1.5 5398.954141141141u,0 5399.930681181181u,0 5399.931681181181u,1.5 5600.326389389389u,1.5 5600.327389389389u,0 5601.303929429429u,0 5601.30492942943u,1.5 5605.21408958959u,1.5 5605.21508958959u,0 5608.146709709709u,0 5608.1477097097095u,1.5 5609.12424974975u,1.5 5609.12524974975u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5664.8440320320315u,1.5 5664.845032032032u,0 5665.821572072072u,0 5665.822572072072u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 5788.991617117117u,1.5 5788.992617117117u,0 5789.9691571571575u,0 5789.970157157158u,1.5 5790.946697197197u,1.5 5790.947697197197u,0 5792.901777277278u,0 5792.902777277278u,1.5 5793.879317317317u,1.5 5793.880317317317u,0 5837.868619119119u,0 5837.869619119119u,1.5 5838.8461591591595u,1.5 5838.84715915916u,0 5840.801239239238u,0 5840.802239239239u,1.5 5888.700701201201u,1.5 5888.701701201201u,0 5889.67824124124u,0 5889.679241241241u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5899.453641641641u,0 5899.4546416416415u,1.5 5900.431181681682u,1.5 5900.432181681682u,0 6101.80442992993u,0 6101.80542992993u,1.5 6102.78196996997u,1.5 6102.7829699699705u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6106.69213013013u,0 6106.69313013013u,1.5 6107.66967017017u,1.5 6107.6706701701705u,0 6108.64721021021u,0 6108.64821021021u,1.5 6159.4792922922925u,1.5 6159.480292292293u,0 6160.456832332332u,0 6160.457832332332u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6208.3562942942945u,0 6208.357294294295u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6291.447197697697u,0 6291.448197697698u,1.5 6337.391579579579u,1.5 6337.392579579579u,0 6339.34665965966u,0 6339.34765965966u,1.5 6340.324199699699u,1.5 6340.3251996997u,0 6342.27927977978u,0 6342.28027977978u,1.5 6343.25681981982u,1.5 6343.25781981982u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6397.021522022022u,0 6397.022522022022u,1.5 6600.34985035035u,1.5 6600.35085035035u,0 6601.32739039039u,0 6601.32839039039u,1.5 6604.26001051051u,1.5 6604.2610105105105u,0 6606.215090590591u,0 6606.216090590591u,1.5 6607.19263063063u,1.5 6607.193630630631u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6664.867492992993u,1.5 6664.868492992993u,0 6665.845033033032u,0 6665.846033033033u,1.5 6705.924174674675u,1.5 6705.925174674675u,0 6706.901714714714u,0 6706.902714714714u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6708.856794794795u,0 6708.857794794795u,1.5 6709.834334834834u,1.5 6709.835334834835u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6752.846096596597u,0 6752.847096596597u,1.5 6791.947698198198u,1.5 6791.948698198198u,0 6835.937u,0 6835.938u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6839.8471601601605u,0 6839.848160160161u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6893.611862362362u,0 6893.612862362363u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0
vb15 b15 0 pwl 0,0  158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 164.22622672672674u,0 164.2272267267267u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 335.2957337337337u,0 335.2967337337337u,1.5 336.2732737737738u,1.5 336.27427377377376u,0 337.2508138138138u,0 337.2518138138138u,1.5 338.2283538538539u,1.5 338.22935385385387u,0 340.18343393393394u,0 340.1844339339339u,1.5 660.816567067067u,1.5 660.817567067067u,0 661.7941071071072u,0 661.7951071071071u,1.5 662.7716471471472u,1.5 662.7726471471472u,0 663.7491871871872u,0 663.7501871871872u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 841.6614744744745u,1.5 841.6624744744745u,0 1161.3170675675676u,0 1161.3180675675678u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1163.2721476476477u,0 1163.2731476476479u,1.5 1164.2496876876876u,1.5 1164.2506876876878u,0 1165.2272277277275u,0 1165.2282277277277u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1254.1833713713713u,1.5 1254.1843713713715u,0 1338.251814814815u,0 1338.252814814815u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1342.1619749749748u,0 1342.162974974975u,1.5 1662.795108108108u,1.5 1662.7961081081082u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1752.7287917917918u,0 1752.729791791792u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1839.7298553553553u,1.5 1839.7308553553555u,0 2162.3180685685684u,0 2162.3190685685686u,1.5 2163.2956086086083u,1.5 2163.2966086086085u,0 2164.2731486486487u,0 2164.274148648649u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2254.2068323323324u,1.5 2254.2078323323326u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2340.2303558558556u,1.5 2340.231355855856u,0 2341.207895895896u,0 2341.208895895896u,1.5 2657.9308688688684u,1.5 2657.9318688688686u,0 2658.9084089089088u,0 2658.909408908909u,1.5 2659.8859489489487u,1.5 2659.886948948949u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2665.751189189189u,0 2665.7521891891893u,1.5 2666.7287292292294u,1.5 2666.7297292292296u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2750.7971726726723u,0 2750.7981726726725u,1.5 2751.7747127127127u,1.5 2751.775712712713u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2839.753316316316u,0 2839.7543163163164u,1.5 2840.730856356356u,1.5 2840.7318563563563u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3335.366116616616u,0 3335.3671166166164u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3836.844157157157u,0 3836.8451571571572u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 4161.38745045045u,0 4161.38845045045u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4336.367117617618u,0 4336.368117617618u,1.5 4337.344657657658u,1.5 4337.345657657658u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4342.232357857858u,0 4342.233357857858u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4840.777778278279u,0 4840.778778278279u,1.5 4841.755318318318u,1.5 4841.756318318318u,0 5160.433371371371u,0 5160.4343713713715u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5162.388451451451u,0 5162.389451451451u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5337.368118618619u,0 5337.369118618619u,1.5 5338.345658658659u,1.5 5338.346658658659u,0 5339.323198698698u,0 5339.324198698699u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5664.8440320320315u,0 5664.845032032032u,1.5 5665.821572072072u,1.5 5665.822572072072u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5838.8461591591595u,0 5838.84715915916u,1.5 5840.801239239238u,1.5 5840.802239239239u,0 6159.4792922922925u,0 6159.480292292293u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6162.411912412412u,0 6162.412912412412u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6337.391579579579u,0 6337.392579579579u,1.5 6339.34665965966u,1.5 6339.34765965966u,0 6340.324199699699u,0 6340.3251996997u,1.5 6342.27927977978u,1.5 6342.28027977978u,0 6343.25681981982u,0 6343.25781981982u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6664.867492992993u,0 6664.868492992993u,1.5 6665.845033033032u,1.5 6665.846033033033u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6752.846096596597u,0 6752.847096596597u,1.5 6835.937u,1.5 6835.938u,0 6837.89208008008u,0 6837.89308008008u,1.5 6839.8471601601605u,1.5 6839.848160160161u,0
vb16 b16 0 pwl 0,0  249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1254.1833713713713u,0 1254.1843713713715u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1752.7287917917918u,1.5 1752.729791791792u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2254.2068323323324u,0 2254.2078323323326u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2750.7971726726723u,1.5 2750.7981726726725u,0 2751.7747127127127u,0 2751.775712712713u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 4251.321134134134u,0 4251.322134134134u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 5250.367055055054u,0 5250.368055055054u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6752.846096596597u,1.5 6752.847096596597u,0

vbb11 bb11 0 pwl 0,1.5  0.9770400400400401u,1.5 0.97804004004004u,0 1.95458008008008u,0 1.95558008008008u,1.5 2.93212012012012u,1.5 2.9331201201201202u,0 3.90966016016016u,0 3.9106601601601603u,1.5 4.8872002002002u,1.5 4.8882002002002u,0 9.7749004004004u,0 9.7759004004004u,1.5 11.72998048048048u,1.5 11.730980480480481u,0 12.70752052052052u,0 12.708520520520521u,1.5 13.68506056056056u,1.5 13.686060560560561u,0 17.59522072072072u,0 17.59622072072072u,1.5 18.572760760760765u,1.5 18.573760760760763u,0 25.415541041041042u,0 25.41654104104104u,1.5 26.393081081081085u,1.5 26.394081081081083u,0 27.370621121121122u,0 27.37162112112112u,1.5 28.348161161161162u,1.5 28.34916116116116u,0 30.303241241241246u,0 30.304241241241243u,1.5 31.280781281281282u,1.5 31.28178128128128u,0 33.23586136136136u,0 33.23686136136136u,1.5 35.19094144144144u,1.5 35.19194144144144u,0 36.16848148148148u,0 36.16948148148148u,1.5 37.146021521521526u,1.5 37.14702152152153u,0 39.1011016016016u,0 39.1021016016016u,1.5 40.07864164164164u,1.5 40.07964164164164u,0 42.03372172172172u,0 42.03472172172172u,1.5 44.966341841841846u,1.5 44.96734184184185u,0 45.94388188188188u,0 45.944881881881884u,1.5 47.89896196196196u,1.5 47.899961961961964u,0 48.876502002002u,0 48.877502002002004u,1.5 50.83158208208208u,1.5 50.832582082082084u,0 52.786662162162166u,0 52.78766216216217u,1.5 53.7642022022022u,1.5 53.765202202202204u,0 54.74174224224224u,0 54.742742242242244u,1.5 55.71928228228228u,1.5 55.720282282282284u,0 58.6519024024024u,0 58.652902402402404u,1.5 59.62944244244244u,1.5 59.630442442442444u,0 63.539602602602606u,0 63.54060260260261u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 71.35992292292292u,1.5 71.36092292292292u,0 72.33746296296296u,0 72.33846296296296u,1.5 76.24762312312312u,1.5 76.24862312312312u,0 78.2027032032032u,0 78.2037032032032u,1.5 80.15778328328328u,1.5 80.15878328328328u,0 85.04548348348348u,0 85.04648348348348u,1.5 86.02302352352352u,1.5 86.02402352352352u,0 87.00056356356356u,0 87.00156356356356u,1.5 90.91072372372372u,1.5 90.91172372372372u,0 92.8658038038038u,0 92.8668038038038u,1.5 94.82088388388388u,1.5 94.82188388388388u,0 95.79842392392392u,0 95.79942392392392u,1.5 96.77596396396396u,1.5 96.77696396396396u,0 97.753504004004u,0 97.754504004004u,1.5 98.73104404404404u,1.5 98.73204404404404u,0 100.68612412412412u,0 100.68712412412413u,1.5 101.66366416416416u,1.5 101.66466416416417u,0 104.59628428428428u,0 104.59728428428429u,1.5 106.55136436436436u,1.5 106.55236436436437u,0 107.5289044044044u,0 107.5299044044044u,1.5 109.48398448448448u,1.5 109.48498448448449u,0 111.43906456456456u,0 111.44006456456457u,1.5 114.37168468468468u,1.5 114.37268468468469u,0 115.34922472472472u,0 115.35022472472473u,1.5 117.3043048048048u,1.5 117.3053048048048u,0 123.16954504504503u,0 123.17054504504503u,1.5 124.14708508508508u,1.5 124.14808508508509u,0 125.12462512512512u,0 125.12562512512513u,1.5 127.07970520520522u,1.5 127.08070520520522u,0 128.05724524524524u,0 128.05824524524522u,1.5 130.01232532532532u,1.5 130.0133253253253u,0 135.8775655655656u,0 135.87856556556557u,1.5 136.85510560560562u,1.5 136.8561056056056u,0 137.83264564564567u,0 137.83364564564565u,1.5 139.78772572572572u,1.5 139.7887257257257u,0 140.76526576576578u,0 140.76626576576575u,1.5 141.74280580580583u,1.5 141.7438058058058u,0 142.72034584584586u,0 142.72134584584583u,1.5 143.69788588588588u,1.5 143.69888588588586u,0 144.67542592592594u,0 144.6764259259259u,1.5 145.65296596596596u,1.5 145.65396596596594u,0 150.54066616616618u,0 150.54166616616615u,1.5 152.49574624624626u,1.5 152.49674624624623u,0 153.4732862862863u,0 153.4742862862863u,1.5 156.40590640640642u,1.5 156.4069064064064u,0 158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 165.20376676676676u,0 165.20476676676674u,1.5 168.1363868868869u,1.5 168.13738688688687u,0 169.11392692692695u,0 169.11492692692693u,1.5 170.09146696696698u,1.5 170.09246696696695u,0 174.97916716716716u,0 174.98016716716714u,1.5 178.88932732732735u,1.5 178.89032732732733u,0 184.7545675675676u,0 184.75556756756757u,1.5 185.73210760760762u,1.5 185.7331076076076u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 189.64226776776778u,0 189.64326776776775u,1.5 190.6198078078078u,1.5 190.62080780780778u,0 191.59734784784786u,0 191.59834784784783u,1.5 192.57488788788788u,1.5 192.57588788788786u,0 194.529967967968u,0 194.53096796796797u,1.5 197.4625880880881u,1.5 197.46358808808807u,0 198.44012812812815u,0 198.44112812812813u,1.5 201.37274824824826u,1.5 201.37374824824823u,0 203.32782832832834u,0 203.3288283283283u,1.5 204.3053683683684u,1.5 204.30636836836837u,0 207.2379884884885u,0 207.23898848848847u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 210.17060860860863u,0 210.1716086086086u,1.5 211.1481486486487u,1.5 211.14914864864866u,0 212.12568868868868u,0 212.12668868868866u,1.5 214.0807687687688u,1.5 214.08176876876877u,0 218.96846896896898u,0 218.96946896896895u,1.5 219.94600900900903u,1.5 219.947009009009u,0 220.92354904904906u,0 220.92454904904903u,1.5 223.85616916916916u,1.5 223.85716916916914u,0 229.72140940940943u,0 229.7224094094094u,1.5 230.69894944944946u,1.5 230.69994944944943u,0 231.6764894894895u,0 231.6774894894895u,1.5 233.63156956956956u,1.5 233.63256956956954u,0 234.60910960960962u,0 234.6101096096096u,1.5 236.5641896896897u,1.5 236.56518968968967u,0 237.54172972972972u,0 237.5427297297297u,1.5 238.51926976976978u,1.5 238.52026976976975u,0 239.4968098098098u,0 239.49780980980978u,1.5 240.47434984984986u,1.5 240.47534984984983u,0 241.4518898898899u,0 241.4528898898899u,1.5 242.42942992992997u,1.5 242.43042992992994u,0 243.40696996996996u,0 243.40796996996994u,1.5 245.36205005005007u,1.5 245.36305005005005u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 256.11499049049047u,1.5 256.11599049049045u,0 259.04761061061066u,0 259.04861061061064u,1.5 260.02515065065063u,1.5 260.0261506506506u,0 261.00269069069066u,0 261.00369069069063u,1.5 261.98023073073074u,1.5 261.9812307307307u,0 263.93531081081085u,0 263.9363108108108u,1.5 265.8903908908909u,1.5 265.8913908908909u,0 270.77809109109114u,0 270.7790910910911u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 272.73317117117114u,0 272.7341711711711u,1.5 275.6657912912913u,1.5 275.6667912912913u,0 279.57595145145143u,0 279.5769514514514u,1.5 280.5534914914915u,1.5 280.5544914914915u,0 281.53103153153154u,0 281.5320315315315u,1.5 282.50857157157157u,1.5 282.50957157157154u,0 283.48611161161165u,0 283.4871116116116u,1.5 287.39627177177175u,1.5 287.3972717717717u,0 289.35135185185186u,0 289.35235185185184u,1.5 290.32889189189194u,1.5 290.3298918918919u,0 294.23905205205205u,0 294.240052052052u,1.5 297.17167217217224u,1.5 297.1726721721722u,0 298.1492122122122u,0 298.1502122122122u,1.5 300.1042922922923u,1.5 300.1052922922923u,0 302.0593723723724u,0 302.0603723723724u,1.5 304.0144524524524u,1.5 304.0154524524524u,0 307.92461261261263u,0 307.9256126126126u,1.5 308.90215265265266u,1.5 308.90315265265264u,0 313.78985285285285u,0 313.7908528528528u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 315.74493293293295u,0 315.74593293293293u,1.5 317.700013013013u,1.5 317.701013013013u,0 318.67755305305303u,0 318.678553053053u,1.5 320.63263313313314u,1.5 320.6336331331331u,0 321.6101731731732u,0 321.6111731731732u,1.5 322.5877132132132u,1.5 322.58871321321317u,0 323.5652532532532u,0 323.5662532532532u,1.5 324.5427932932933u,1.5 324.5437932932933u,0 326.4978733733734u,0 326.4988733733734u,1.5 328.45295345345346u,1.5 328.45395345345344u,0 330.4080335335335u,0 330.4090335335335u,1.5 332.3631136136136u,1.5 332.3641136136136u,0 333.3406536536537u,0 333.3416536536537u,1.5 334.31819369369373u,1.5 334.3191936936937u,0 335.2957337337337u,0 335.2967337337337u,1.5 336.2732737737738u,1.5 336.27427377377376u,0 337.2508138138138u,0 337.2518138138138u,1.5 338.2283538538539u,1.5 338.22935385385387u,0 340.18343393393394u,0 340.1844339339339u,1.5 343.1160540540541u,1.5 343.11705405405405u,0 344.0935940940941u,0 344.0945940940941u,1.5 345.0711341341341u,1.5 345.0721341341341u,0 349.9588343343343u,0 349.9598343343343u,1.5 350.9363743743744u,1.5 350.9373743743744u,0 353.8689944944945u,0 353.86999449449445u,1.5 354.8465345345345u,1.5 354.8475345345345u,0 355.8240745745746u,0 355.82507457457456u,1.5 357.7791546546547u,1.5 357.78015465465467u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 367.55455505505506u,1.5 367.55555505505504u,0 368.5320950950951u,0 368.53309509509506u,1.5 371.4647152152152u,1.5 371.4657152152152u,0 372.44225525525525u,0 372.4432552552552u,1.5 375.3748753753754u,1.5 375.37587537537536u,0 378.3074954954955u,0 378.3084954954955u,1.5 380.26257557557557u,1.5 380.26357557557554u,0 381.2401156156156u,0 381.24111561561557u,1.5 386.1278158158158u,1.5 386.12881581581576u,0 388.0828958958959u,0 388.08389589589586u,1.5 390.037975975976u,1.5 390.038975975976u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 395.90321621621626u,0 395.90421621621624u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 398.83583633633634u,0 398.8368363363363u,1.5 399.81337637637637u,1.5 399.81437637637634u,0 400.79091641641645u,0 400.7919164164164u,1.5 401.7684564564565u,1.5 401.76945645645645u,0 402.7459964964965u,0 402.7469964964965u,1.5 403.7235365365366u,1.5 403.72453653653656u,0 404.70107657657655u,0 404.70207657657653u,1.5 406.65615665665666u,1.5 406.65715665665664u,0 407.6336966966967u,0 407.63469669669666u,1.5 409.5887767767768u,1.5 409.5897767767768u,0 410.5663168168168u,0 410.5673168168168u,1.5 411.54385685685685u,1.5 411.5448568568568u,0 412.5213968968969u,0 412.52239689689685u,1.5 414.476476976977u,1.5 414.47747697697696u,0 415.45401701701707u,0 415.45501701701704u,1.5 417.40909709709706u,1.5 417.41009709709704u,0 418.38663713713714u,0 418.3876371371371u,1.5 422.29679729729736u,1.5 422.29779729729734u,0 424.25187737737735u,0 424.25287737737733u,1.5 425.22941741741744u,1.5 425.2304174174174u,0 427.18449749749755u,0 427.1854974974975u,1.5 428.16203753753757u,1.5 428.16303753753755u,0 432.07219769769773u,0 432.0731976976977u,1.5 433.04973773773776u,1.5 433.05073773773773u,0 434.0272777777778u,0 434.02827777777776u,1.5 435.00481781781787u,1.5 435.00581781781784u,0 435.98235785785783u,0 435.9833578578578u,1.5 437.93743793793794u,1.5 437.9384379379379u,0 438.91497797797797u,0 438.91597797797795u,1.5 449.6679184184184u,1.5 449.6689184184184u,0 450.64545845845845u,0 450.6464584584584u,1.5 451.62299849849853u,1.5 451.6239984984985u,0 452.60053853853856u,0 452.60153853853853u,1.5 453.5780785785786u,1.5 453.57907857857856u,0 455.53315865865864u,0 455.5341586586586u,1.5 456.5106986986987u,1.5 456.5116986986987u,0 460.4208588588588u,0 460.4218588588588u,1.5 461.3983988988989u,1.5 461.3993988988989u,0 462.37593893893893u,0 462.3769389389389u,1.5 463.353478978979u,1.5 463.354478978979u,0 466.28609909909915u,0 466.2870990990991u,1.5 468.2411791791792u,1.5 468.2421791791792u,0 470.19625925925925u,0 470.1972592592592u,1.5 471.17379929929933u,1.5 471.1747992992993u,0 472.15133933933936u,0 472.15233933933933u,1.5 474.1064194194194u,1.5 474.1074194194194u,0 475.08395945945944u,0 475.0849594594594u,1.5 476.0614994994995u,1.5 476.0624994994995u,0 478.0165795795796u,0 478.0175795795796u,1.5 484.8593598598599u,1.5 484.8603598598599u,0 485.8368998998999u,0 485.83789989989987u,1.5 486.8144399399399u,1.5 486.8154399399399u,0 487.79197997998u,0 487.79297997998u,1.5 488.7695200200201u,1.5 488.77052002002006u,0 489.7470600600601u,0 489.7480600600601u,1.5 495.6123003003003u,1.5 495.6133003003003u,0 497.56738038038037u,0 497.56838038038035u,1.5 499.5224604604605u,1.5 499.52346046046046u,0 500.5000005005005u,0 500.5010005005005u,1.5 503.4326206206207u,1.5 503.4336206206207u,0 504.41016066066067u,0 504.41116066066064u,1.5 507.34278078078074u,1.5 507.3437807807807u,0 508.3203208208209u,0 508.32132082082086u,1.5 509.2978608608609u,1.5 509.2988608608609u,0 510.2754009009009u,0 510.27640090090085u,1.5 518.0957212212213u,1.5 518.0967212212213u,0 519.0732612612613u,0 519.0742612612613u,1.5 521.0283413413413u,1.5 521.0293413413413u,0 522.0058813813813u,0 522.0068813813813u,1.5 525.9160415415415u,1.5 525.9170415415415u,0 526.8935815815815u,0 526.8945815815815u,1.5 528.8486616616617u,1.5 528.8496616616617u,0 530.8037417417418u,0 530.8047417417417u,1.5 531.7812817817818u,1.5 531.7822817817818u,0 533.7363618618618u,0 533.7373618618618u,1.5 534.7139019019019u,1.5 534.7149019019018u,0 540.5791421421421u,0 540.5801421421421u,1.5 542.5342222222223u,1.5 542.5352222222223u,0 545.4668423423423u,0 545.4678423423422u,1.5 546.4443823823824u,1.5 546.4453823823824u,0 547.4219224224224u,0 547.4229224224224u,1.5 548.3994624624625u,1.5 548.4004624624624u,0 549.3770025025025u,0 549.3780025025025u,1.5 550.3545425425425u,1.5 550.3555425425425u,0 551.3320825825826u,0 551.3330825825826u,1.5 553.2871626626627u,1.5 553.2881626626627u,0 554.2647027027027u,0 554.2657027027027u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 561.107482982983u,0 561.108482982983u,1.5 563.0625630630631u,1.5 563.063563063063u,0 564.0401031031031u,0 564.0411031031031u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 568.9278033033033u,0 568.9288033033033u,1.5 569.9053433433434u,1.5 569.9063433433433u,0 575.7705835835836u,0 575.7715835835836u,1.5 576.7481236236237u,1.5 576.7491236236236u,0 577.7256636636637u,0 577.7266636636637u,1.5 584.5684439439439u,1.5 584.5694439439438u,0 585.545983983984u,0 585.546983983984u,1.5 587.501064064064u,1.5 587.502064064064u,0 589.4561441441441u,0 589.4571441441441u,1.5 590.4336841841842u,1.5 590.4346841841842u,0 592.3887642642643u,0 592.3897642642643u,1.5 594.3438443443445u,1.5 594.3448443443444u,0 595.3213843843844u,0 595.3223843843843u,1.5 598.2540045045045u,1.5 598.2550045045044u,0 599.2315445445446u,0 599.2325445445446u,1.5 600.2090845845846u,1.5 600.2100845845846u,0 601.1866246246246u,0 601.1876246246246u,1.5 602.1641646646647u,1.5 602.1651646646646u,0 603.1417047047047u,0 603.1427047047047u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 606.0743248248249u,0 606.0753248248249u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 613.8946451451452u,0 613.8956451451452u,1.5 615.8497252252253u,1.5 615.8507252252252u,0 616.8272652652653u,0 616.8282652652653u,1.5 620.7374254254254u,1.5 620.7384254254254u,0 621.7149654654654u,0 621.7159654654654u,1.5 623.6700455455456u,1.5 623.6710455455456u,0 628.5577457457458u,0 628.5587457457458u,1.5 637.355606106106u,1.5 637.356606106106u,0 643.2208463463464u,0 643.2218463463464u,1.5 645.1759264264264u,1.5 645.1769264264263u,0 646.1534664664664u,0 646.1544664664664u,1.5 649.0860865865866u,1.5 649.0870865865866u,0 653.9737867867868u,0 653.9747867867868u,1.5 654.9513268268269u,1.5 654.9523268268268u,0 656.9064069069069u,0 656.9074069069069u,1.5 660.816567067067u,1.5 660.817567067067u,0 661.7941071071072u,0 661.7951071071071u,1.5 662.7716471471472u,1.5 662.7726471471472u,0 663.7491871871872u,0 663.7501871871872u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 666.6818073073074u,0 666.6828073073074u,1.5 667.6593473473474u,1.5 667.6603473473474u,0 670.5919674674674u,0 670.5929674674674u,1.5 672.5470475475475u,1.5 672.5480475475475u,0 674.5021276276276u,0 674.5031276276276u,1.5 675.4796676676676u,1.5 675.4806676676676u,0 678.4122877877878u,0 678.4132877877878u,1.5 679.3898278278278u,1.5 679.3908278278278u,0 680.3673678678679u,0 680.3683678678678u,1.5 682.3224479479479u,1.5 682.3234479479479u,0 683.299987987988u,0 683.3009879879879u,1.5 685.255068068068u,1.5 685.256068068068u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 692.0978483483484u,0 692.0988483483484u,1.5 696.0080085085085u,1.5 696.0090085085085u,0 696.9855485485485u,0 696.9865485485485u,1.5 697.9630885885886u,1.5 697.9640885885885u,0 703.8283288288288u,0 703.8293288288288u,1.5 707.7384889889889u,1.5 707.7394889889889u,0 708.716029029029u,0 708.7170290290289u,1.5 709.693569069069u,1.5 709.694569069069u,0 712.6261891891892u,0 712.6271891891892u,1.5 713.6037292292292u,1.5 713.6047292292292u,0 714.5812692692692u,0 714.5822692692692u,1.5 716.5363493493494u,1.5 716.5373493493494u,0 717.5138893893894u,0 717.5148893893894u,1.5 718.4914294294294u,1.5 718.4924294294294u,0 722.4015895895895u,0 722.4025895895895u,1.5 723.3791296296296u,1.5 723.3801296296296u,0 724.3566696696697u,0 724.3576696696697u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 729.24436986987u,1.5 729.2453698698699u,0 730.22190990991u,0 730.22290990991u,1.5 731.19944994995u,1.5 731.20044994995u,0 733.15453003003u,0 733.1555300300299u,1.5 734.1320700700701u,1.5 734.1330700700701u,0 735.1096101101101u,0 735.1106101101101u,1.5 736.0871501501501u,1.5 736.0881501501501u,0 737.0646901901902u,0 737.0656901901901u,1.5 739.0197702702703u,1.5 739.0207702702703u,0 740.9748503503504u,0 740.9758503503504u,1.5 742.9299304304304u,1.5 742.9309304304304u,0 744.8850105105105u,0 744.8860105105105u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 755.637950950951u,0 755.638950950951u,1.5 756.615490990991u,1.5 756.616490990991u,0 757.593031031031u,0 757.594031031031u,1.5 764.4358113113113u,1.5 764.4368113113113u,0 765.4133513513514u,0 765.4143513513513u,1.5 766.3908913913914u,1.5 766.3918913913914u,0 767.3684314314314u,0 767.3694314314314u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 771.2785915915915u,0 771.2795915915915u,1.5 772.2561316316315u,1.5 772.2571316316315u,0 775.1887517517517u,0 775.1897517517517u,1.5 776.1662917917918u,1.5 776.1672917917917u,0 777.1438318318318u,0 777.1448318318318u,1.5 781.053991991992u,1.5 781.054991991992u,0 782.031532032032u,0 782.032532032032u,1.5 783.0090720720721u,1.5 783.010072072072u,0 784.9641521521521u,0 784.9651521521521u,1.5 785.9416921921921u,1.5 785.9426921921921u,0 787.8967722722723u,0 787.8977722722723u,1.5 790.8293923923924u,1.5 790.8303923923924u,0 792.7844724724725u,0 792.7854724724725u,1.5 793.7620125125126u,1.5 793.7630125125125u,0 796.6946326326326u,0 796.6956326326326u,1.5 797.6721726726727u,1.5 797.6731726726726u,0 799.6272527527527u,0 799.6282527527527u,1.5 803.5374129129129u,1.5 803.5384129129129u,0 806.4700330330331u,0 806.4710330330331u,1.5 807.4475730730732u,1.5 807.4485730730731u,0 808.4251131131131u,0 808.426113113113u,1.5 814.2903533533533u,1.5 814.2913533533533u,0 815.2678933933934u,0 815.2688933933933u,1.5 817.2229734734735u,1.5 817.2239734734735u,0 821.1331336336336u,0 821.1341336336336u,1.5 824.0657537537537u,1.5 824.0667537537537u,0 832.8636141141141u,0 832.864614114114u,1.5 835.7962342342342u,1.5 835.7972342342342u,0 836.7737742742743u,0 836.7747742742743u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 842.6390145145145u,1.5 842.6400145145145u,0 843.6165545545546u,0 843.6175545545545u,1.5 846.5491746746746u,1.5 846.5501746746746u,0 847.5267147147147u,0 847.5277147147146u,1.5 848.5042547547547u,1.5 848.5052547547547u,0 849.4817947947948u,0 849.4827947947948u,1.5 851.4368748748749u,1.5 851.4378748748749u,0 852.4144149149149u,0 852.4154149149149u,1.5 853.3919549549549u,1.5 853.3929549549549u,0 854.3694949949951u,0 854.370494994995u,1.5 859.2571951951952u,1.5 859.2581951951952u,0 860.2347352352352u,0 860.2357352352352u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 868.0550555555556u,0 868.0560555555555u,1.5 870.0101356356357u,1.5 870.0111356356357u,0 870.9876756756756u,0 870.9886756756756u,1.5 878.8079959959961u,1.5 878.808995995996u,0 882.7181561561562u,0 882.7191561561561u,1.5 883.6956961961962u,1.5 883.6966961961962u,0 886.6283163163163u,0 886.6293163163162u,1.5 894.4486366366367u,1.5 894.4496366366367u,0 896.4037167167166u,0 896.4047167167166u,1.5 897.3812567567567u,1.5 897.3822567567566u,0 902.2689569569569u,0 902.2699569569569u,1.5 904.2240370370371u,1.5 904.225037037037u,0 905.2015770770771u,0 905.2025770770771u,1.5 907.1566571571572u,1.5 907.1576571571571u,0 909.1117372372372u,0 909.1127372372372u,1.5 911.0668173173173u,1.5 911.0678173173172u,0 912.0443573573574u,0 912.0453573573574u,1.5 913.0218973973974u,1.5 913.0228973973974u,0 913.9994374374375u,0 914.0004374374374u,1.5 915.9545175175175u,1.5 915.9555175175175u,0 916.9320575575576u,0 916.9330575575576u,1.5 917.9095975975977u,1.5 917.9105975975976u,0 919.8646776776777u,0 919.8656776776777u,1.5 921.8197577577578u,1.5 921.8207577577577u,0 923.7748378378378u,0 923.7758378378378u,1.5 924.7523778778778u,1.5 924.7533778778778u,0 925.7299179179179u,0 925.7309179179178u,1.5 927.684997997998u,1.5 927.685997997998u,0 928.6625380380381u,0 928.663538038038u,1.5 932.5726981981983u,1.5 932.5736981981983u,0 933.5502382382382u,0 933.5512382382382u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 938.4379384384384u,0 938.4389384384384u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 947.2357987987988u,0 947.2367987987988u,1.5 948.2133388388388u,1.5 948.2143388388388u,0 949.1908788788788u,0 949.1918788788788u,1.5 950.1684189189189u,1.5 950.1694189189188u,0 951.145958958959u,0 951.146958958959u,1.5 957.0111991991993u,1.5 957.0121991991992u,0 957.9887392392392u,0 957.9897392392392u,1.5 959.9438193193192u,1.5 959.9448193193192u,0 960.9213593593594u,0 960.9223593593593u,1.5 964.8315195195195u,1.5 964.8325195195195u,0 966.7865995995996u,0 966.7875995995996u,1.5 967.7641396396397u,1.5 967.7651396396396u,0 968.7416796796797u,0 968.7426796796797u,1.5 970.6967597597597u,1.5 970.6977597597597u,0 972.6518398398398u,0 972.6528398398398u,1.5 973.6293798798798u,1.5 973.6303798798798u,0 974.60691991992u,0 974.6079199199199u,1.5 975.58445995996u,1.5 975.58545995996u,0 977.5395400400402u,0 977.5405400400401u,1.5 978.5170800800801u,1.5 978.51808008008u,0 981.4497002002003u,0 981.4507002002002u,1.5 984.3823203203203u,1.5 984.3833203203203u,0 986.3374004004004u,0 986.3384004004004u,1.5 987.3149404404405u,1.5 987.3159404404405u,0 989.2700205205206u,0 989.2710205205206u,1.5 992.2026406406408u,1.5 992.2036406406407u,0 993.1801806806807u,0 993.1811806806807u,1.5 995.1352607607607u,1.5 995.1362607607607u,0 999.045420920921u,0 999.0464209209209u,1.5 1000.0229609609609u,1.5 1000.0239609609608u,0 1001.9780410410411u,0 1001.9790410410411u,1.5 1002.955581081081u,1.5 1002.956581081081u,0 1003.9331211211212u,0 1003.9341211211212u,1.5 1005.8882012012012u,1.5 1005.8892012012012u,0 1006.8657412412414u,0 1006.8667412412414u,1.5 1007.8432812812813u,1.5 1007.8442812812813u,0 1013.7085215215216u,0 1013.7095215215215u,1.5 1014.6860615615615u,1.5 1014.6870615615614u,0 1016.6411416416418u,0 1016.6421416416417u,1.5 1017.6186816816817u,1.5 1017.6196816816816u,0 1021.5288418418419u,0 1021.5298418418419u,1.5 1022.5063818818818u,1.5 1022.5073818818818u,0 1026.416542042042u,0 1026.4175420420422u,1.5 1027.394082082082u,1.5 1027.3950820820821u,0 1028.371622122122u,0 1028.3726221221223u,1.5 1029.349162162162u,1.5 1029.3501621621622u,0 1030.3267022022021u,0 1030.3277022022023u,1.5 1031.3042422422423u,1.5 1031.3052422422425u,0 1032.2817822822822u,0 1032.2827822822824u,1.5 1033.2593223223223u,1.5 1033.2603223223225u,0 1034.2368623623622u,0 1034.2378623623624u,1.5 1041.0796426426425u,1.5 1041.0806426426427u,0 1042.0571826826824u,0 1042.0581826826826u,1.5 1045.9673428428428u,1.5 1045.968342842843u,0 1046.9448828828827u,0 1046.9458828828829u,1.5 1047.9224229229228u,1.5 1047.923422922923u,0 1048.8999629629627u,0 1048.900962962963u,1.5 1049.8775030030029u,1.5 1049.878503003003u,0 1050.855043043043u,0 1050.8560430430432u,1.5 1051.832583083083u,1.5 1051.833583083083u,0 1052.810123123123u,0 1052.8111231231233u,1.5 1053.787663163163u,1.5 1053.7886631631632u,0 1054.765203203203u,0 1054.7662032032033u,1.5 1055.7427432432432u,1.5 1055.7437432432434u,0 1057.6978233233233u,0 1057.6988233233235u,1.5 1058.6753633633632u,1.5 1058.6763633633634u,0 1061.6079834834834u,0 1061.6089834834836u,1.5 1062.5855235235235u,1.5 1062.5865235235237u,0 1065.5181436436435u,0 1065.5191436436437u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1070.4058438438437u,1.5 1070.406843843844u,0 1071.3833838838837u,0 1071.3843838838839u,1.5 1077.248624124124u,1.5 1077.2496241241242u,0 1079.203704204204u,0 1079.2047042042043u,1.5 1080.1812442442442u,1.5 1080.1822442442444u,0 1081.1587842842841u,0 1081.1597842842843u,1.5 1082.1363243243243u,1.5 1082.1373243243245u,0 1086.0464844844844u,0 1086.0474844844846u,1.5 1087.0240245245245u,1.5 1087.0250245245247u,0 1093.8668048048046u,0 1093.8678048048048u,1.5 1096.7994249249248u,1.5 1096.800424924925u,0 1102.6646651651652u,0 1102.6656651651654u,1.5 1103.642205205205u,1.5 1103.6432052052053u,0 1104.6197452452452u,0 1104.6207452452454u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1107.5523653653654u,0 1107.5533653653656u,1.5 1108.5299054054053u,1.5 1108.5309054054055u,0 1109.5074454454455u,0 1109.5084454454457u,1.5 1113.4176056056056u,1.5 1113.4186056056058u,0 1115.3726856856854u,0 1115.3736856856856u,1.5 1116.3502257257255u,1.5 1116.3512257257257u,0 1119.2828458458457u,0 1119.283845845846u,1.5 1121.2379259259258u,1.5 1121.238925925926u,0 1122.215465965966u,0 1122.216465965966u,1.5 1124.170546046046u,1.5 1124.1715460460462u,0 1125.1480860860859u,0 1125.149086086086u,1.5 1126.125626126126u,1.5 1126.1266261261262u,0 1127.1031661661661u,0 1127.1041661661664u,1.5 1130.035786286286u,1.5 1130.0367862862863u,0 1131.0133263263263u,0 1131.0143263263265u,1.5 1131.9908663663664u,1.5 1131.9918663663666u,0 1134.9234864864864u,0 1134.9244864864866u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1142.7438068068066u,1.5 1142.7448068068068u,0 1143.7213468468467u,0 1143.722346846847u,1.5 1144.6988868868866u,1.5 1144.6998868868868u,0 1148.609047047047u,0 1148.6100470470471u,1.5 1150.564127127127u,1.5 1150.5651271271272u,0 1156.4293673673674u,0 1156.4303673673676u,1.5 1158.3844474474474u,1.5 1158.3854474474476u,0 1161.3170675675676u,0 1161.3180675675678u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1165.2272277277275u,0 1165.2282277277277u,1.5 1166.2047677677676u,1.5 1166.2057677677678u,0 1167.1823078078075u,0 1167.1833078078078u,1.5 1170.1149279279277u,1.5 1170.115927927928u,0 1172.0700080080078u,0 1172.071008008008u,1.5 1173.047548048048u,1.5 1173.0485480480481u,0 1175.002628128128u,0 1175.0036281281282u,1.5 1176.957708208208u,1.5 1176.9587082082082u,0 1178.912788288288u,0 1178.9137882882883u,1.5 1179.8903283283282u,1.5 1179.8913283283284u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1190.6432687687686u,1.5 1190.6442687687688u,0 1191.6208088088085u,0 1191.6218088088087u,1.5 1192.5983488488487u,1.5 1192.5993488488489u,0 1197.486049049049u,0 1197.4870490490491u,1.5 1199.441129129129u,1.5 1199.4421291291292u,0 1200.418669169169u,0 1200.4196691691693u,1.5 1201.396209209209u,1.5 1201.3972092092092u,0 1202.3737492492492u,0 1202.3747492492494u,1.5 1203.3512892892893u,1.5 1203.3522892892895u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1208.2389894894895u,1.5 1208.2399894894897u,0 1210.1940695695696u,0 1210.1950695695698u,1.5 1213.1266896896898u,1.5 1213.12768968969u,0 1214.1042297297297u,0 1214.10522972973u,1.5 1215.0817697697696u,1.5 1215.0827697697698u,0 1217.0368498498497u,0 1217.0378498498499u,1.5 1218.0143898898898u,1.5 1218.01538988989u,0 1218.9919299299297u,0 1218.99292992993u,1.5 1219.9694699699699u,1.5 1219.97046996997u,0 1220.9470100100098u,0 1220.94801001001u,1.5 1223.87963013013u,1.5 1223.8806301301302u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1232.6774904904905u,0 1232.6784904904907u,1.5 1234.6325705705706u,1.5 1234.6335705705708u,0 1241.4753508508506u,0 1241.4763508508508u,1.5 1242.4528908908908u,1.5 1242.453890890891u,0 1243.4304309309307u,0 1243.431430930931u,1.5 1244.4079709709708u,1.5 1244.408970970971u,0 1245.3855110110107u,0 1245.386511011011u,1.5 1246.363051051051u,1.5 1246.364051051051u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1260.0486116116115u,0 1260.0496116116117u,1.5 1261.0261516516516u,1.5 1261.0271516516518u,0 1262.0036916916918u,0 1262.004691691692u,1.5 1265.9138518518516u,1.5 1265.9148518518518u,0 1266.8913918918918u,0 1266.892391891892u,1.5 1267.8689319319317u,1.5 1267.869931931932u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1271.779092092092u,1.5 1271.7800920920922u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1276.6667922922923u,1.5 1276.6677922922925u,0 1278.6218723723723u,0 1278.6228723723725u,1.5 1279.5994124124122u,1.5 1279.6004124124124u,0 1280.5769524524524u,0 1280.5779524524526u,1.5 1287.4197327327327u,1.5 1287.4207327327329u,0 1288.3972727727728u,0 1288.398272772773u,1.5 1289.3748128128127u,1.5 1289.375812812813u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1291.3298928928928u,1.5 1291.330892892893u,0 1292.3074329329327u,0 1292.3084329329329u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1295.2400530530529u,0 1295.241053053053u,1.5 1298.172673173173u,1.5 1298.1736731731733u,0 1303.0603733733733u,0 1303.0613733733735u,1.5 1305.0154534534533u,1.5 1305.0164534534536u,0 1305.9929934934935u,0 1305.9939934934937u,1.5 1306.9705335335334u,1.5 1306.9715335335336u,0 1307.9480735735735u,0 1307.9490735735737u,1.5 1308.9256136136135u,1.5 1308.9266136136137u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1315.7683938938937u,1.5 1315.769393893894u,0 1316.7459339339337u,0 1316.7469339339339u,1.5 1318.701014014014u,1.5 1318.7020140140141u,0 1319.6785540540538u,0 1319.679554054054u,1.5 1320.656094094094u,1.5 1320.6570940940942u,0 1327.4988743743743u,0 1327.4998743743745u,1.5 1329.4539544544543u,1.5 1329.4549544544545u,0 1332.3865745745745u,0 1332.3875745745747u,1.5 1333.3641146146147u,1.5 1333.3651146146149u,0 1338.251814814815u,0 1338.252814814815u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1343.139515015015u,0 1343.1405150150151u,1.5 1344.1170550550548u,1.5 1344.118055055055u,0 1345.094595095095u,0 1345.0955950950952u,1.5 1346.0721351351349u,1.5 1346.073135135135u,0 1347.049675175175u,0 1347.0506751751752u,1.5 1349.004755255255u,1.5 1349.0057552552553u,0 1350.9598353353351u,0 1350.9608353353353u,1.5 1352.9149154154154u,1.5 1352.9159154154156u,0 1353.8924554554553u,0 1353.8934554554555u,1.5 1356.8250755755755u,1.5 1356.8260755755757u,0 1358.7801556556556u,0 1358.7811556556558u,1.5 1359.7576956956957u,1.5 1359.758695695696u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1367.578016016016u,1.5 1367.579016016016u,0 1368.5555560560558u,0 1368.556556056056u,1.5 1369.533096096096u,1.5 1369.5340960960962u,0 1370.5106361361359u,0 1370.511636136136u,1.5 1371.488176176176u,1.5 1371.4891761761762u,0 1373.443256256256u,0 1373.4442562562563u,1.5 1374.4207962962962u,1.5 1374.4217962962964u,0 1376.3758763763763u,0 1376.3768763763765u,1.5 1377.3534164164164u,1.5 1377.3544164164166u,0 1378.3309564564563u,0 1378.3319564564565u,1.5 1379.3084964964964u,1.5 1379.3094964964966u,0 1380.2860365365364u,0 1380.2870365365366u,1.5 1383.2186566566565u,1.5 1383.2196566566568u,0 1385.1737367367366u,0 1385.1747367367368u,1.5 1386.1512767767767u,1.5 1386.152276776777u,0 1387.1288168168169u,0 1387.129816816817u,1.5 1388.1063568568568u,1.5 1388.107356856857u,0 1392.016517017017u,0 1392.017517017017u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1399.836837337337u,1.5 1399.8378373373373u,0 1403.7469974974974u,0 1403.7479974974976u,1.5 1404.7245375375373u,1.5 1404.7255375375375u,0 1406.6796176176176u,0 1406.6806176176178u,1.5 1407.6571576576575u,1.5 1407.6581576576577u,0 1408.6346976976977u,0 1408.6356976976979u,1.5 1409.6122377377376u,1.5 1409.6132377377378u,0 1411.5673178178179u,0 1411.568317817818u,1.5 1414.4999379379378u,1.5 1414.500937937938u,0 1415.4774779779777u,0 1415.478477977978u,1.5 1418.410098098098u,1.5 1418.4110980980981u,0 1419.3876381381378u,0 1419.388638138138u,1.5 1420.365178178178u,1.5 1420.3661781781782u,0 1421.3427182182181u,0 1421.3437182182183u,1.5 1422.320258258258u,1.5 1422.3212582582582u,0 1423.2977982982982u,0 1423.2987982982984u,1.5 1425.2528783783782u,1.5 1425.2538783783784u,0 1426.2304184184184u,0 1426.2314184184186u,1.5 1427.2079584584583u,1.5 1427.2089584584585u,0 1430.1405785785785u,0 1430.1415785785787u,1.5 1432.0956586586585u,1.5 1432.0966586586587u,0 1433.0731986986987u,0 1433.0741986986989u,1.5 1434.0507387387386u,1.5 1434.0517387387388u,0 1436.0058188188189u,0 1436.006818818819u,1.5 1438.938438938939u,1.5 1438.9394389389392u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1440.8935190190189u,1.5 1440.894519019019u,0 1441.8710590590588u,0 1441.872059059059u,1.5 1444.803679179179u,1.5 1444.8046791791792u,0 1445.781219219219u,0 1445.7822192192193u,1.5 1446.758759259259u,1.5 1446.7597592592592u,0 1447.7362992992992u,0 1447.7372992992994u,1.5 1449.6913793793792u,1.5 1449.6923793793794u,0 1450.6689194194194u,0 1450.6699194194196u,1.5 1451.6464594594593u,1.5 1451.6474594594595u,0 1453.6015395395395u,0 1453.6025395395397u,1.5 1454.5790795795795u,1.5 1454.5800795795797u,0 1464.35447997998u,0 1464.3554799799801u,1.5 1465.3320200200199u,1.5 1465.33302002002u,0 1467.2871001001u,0 1467.2881001001u,1.5 1468.26464014014u,1.5 1468.2656401401402u,0 1470.21972022022u,0 1470.2207202202203u,1.5 1471.19726026026u,1.5 1471.1982602602602u,0 1473.1523403403403u,0 1473.1533403403405u,1.5 1474.1298803803802u,1.5 1474.1308803803804u,0 1476.0849604604603u,0 1476.0859604604605u,1.5 1477.0625005005004u,1.5 1477.0635005005006u,0 1478.0400405405405u,0 1478.0410405405407u,1.5 1480.9726606606605u,1.5 1480.9736606606607u,0 1481.9502007007006u,0 1481.9512007007008u,1.5 1482.9277407407408u,1.5 1482.928740740741u,0 1483.9052807807807u,0 1483.906280780781u,1.5 1489.7705210210208u,1.5 1489.771521021021u,0 1490.7480610610608u,0 1490.749061061061u,1.5 1494.658221221221u,1.5 1494.6592212212213u,0 1495.635761261261u,0 1495.6367612612612u,1.5 1510.2988618618617u,1.5 1510.299861861862u,0 1511.2764019019019u,0 1511.277401901902u,1.5 1513.231481981982u,1.5 1513.2324819819821u,0 1514.209022022022u,0 1514.2100220220223u,1.5 1518.119182182182u,1.5 1518.1201821821821u,0 1519.096722222222u,0 1519.0977222222223u,1.5 1520.074262262262u,1.5 1520.0752622622622u,0 1521.0518023023021u,0 1521.0528023023023u,1.5 1522.0293423423423u,1.5 1522.0303423423425u,0 1523.0068823823822u,0 1523.0078823823824u,1.5 1524.9619624624622u,1.5 1524.9629624624624u,0 1525.9395025025024u,0 1525.9405025025026u,1.5 1526.9170425425425u,1.5 1526.9180425425427u,0 1527.8945825825824u,0 1527.8955825825826u,1.5 1530.8272027027026u,1.5 1530.8282027027028u,0 1531.8047427427427u,0 1531.805742742743u,1.5 1532.7822827827827u,1.5 1532.7832827827829u,0 1542.557683183183u,0 1542.5586831831831u,1.5 1543.535223223223u,1.5 1543.5362232232233u,0 1545.490303303303u,0 1545.4913033033033u,1.5 1546.4678433433432u,1.5 1546.4688433433435u,0 1548.4229234234233u,0 1548.4239234234235u,1.5 1549.4004634634632u,1.5 1549.4014634634634u,0 1550.3780035035034u,0 1550.3790035035036u,1.5 1551.3555435435435u,1.5 1551.3565435435437u,0 1552.3330835835834u,0 1552.3340835835836u,1.5 1553.3106236236235u,1.5 1553.3116236236237u,0 1554.2881636636635u,0 1554.2891636636637u,1.5 1562.108483983984u,1.5 1562.109483983984u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1565.041104104104u,1.5 1565.0421041041043u,0 1566.996184184184u,0 1566.997184184184u,1.5 1567.973724224224u,1.5 1567.9747242242242u,0 1575.7940445445445u,0 1575.7950445445447u,1.5 1576.7715845845844u,1.5 1576.7725845845846u,0 1582.6368248248248u,0 1582.637824824825u,1.5 1583.614364864865u,1.5 1583.6153648648651u,0 1585.569444944945u,0 1585.5704449449452u,1.5 1586.5469849849849u,1.5 1586.547984984985u,0 1587.524525025025u,0 1587.5255250250252u,1.5 1589.479605105105u,1.5 1589.4806051051053u,0 1596.3223853853851u,0 1596.3233853853853u,1.5 1597.2999254254253u,1.5 1597.3009254254255u,0 1598.2774654654654u,0 1598.2784654654656u,1.5 1601.2100855855854u,1.5 1601.2110855855856u,0 1603.1651656656657u,0 1603.1661656656659u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1607.0753258258258u,1.5 1607.076325825826u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1613.918106106106u,0 1613.9191061061063u,1.5 1618.805806306306u,1.5 1618.8068063063063u,0 1619.7833463463462u,0 1619.7843463463464u,1.5 1621.7384264264263u,1.5 1621.7394264264265u,0 1628.5812067067066u,0 1628.5822067067068u,1.5 1629.5587467467467u,1.5 1629.559746746747u,0 1630.5362867867866u,0 1630.5372867867868u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1641.289227227227u,0 1641.2902272272272u,1.5 1642.2667672672671u,1.5 1642.2677672672673u,0 1643.244307307307u,0 1643.2453073073073u,1.5 1644.2218473473472u,1.5 1644.2228473473474u,0 1645.199387387387u,0 1645.2003873873873u,1.5 1650.0870875875873u,1.5 1650.0880875875876u,0 1651.0646276276275u,0 1651.0656276276277u,1.5 1652.0421676676676u,1.5 1652.0431676676678u,0 1654.9747877877876u,0 1654.9757877877878u,1.5 1656.9298678678679u,1.5 1656.930867867868u,0 1657.9074079079078u,0 1657.908407907908u,1.5 1662.795108108108u,1.5 1662.7961081081082u,0 1665.727728228228u,0 1665.7287282282282u,1.5 1666.7052682682681u,1.5 1666.7062682682683u,0 1668.6603483483482u,0 1668.6613483483484u,1.5 1674.5255885885883u,1.5 1674.5265885885885u,0 1675.5031286286285u,0 1675.5041286286287u,1.5 1677.4582087087085u,1.5 1677.4592087087087u,0 1678.4357487487487u,0 1678.4367487487489u,1.5 1679.4132887887886u,1.5 1679.4142887887888u,0 1680.3908288288287u,0 1680.391828828829u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1689.1886891891893u,0 1689.1896891891895u,1.5 1691.1437692692691u,1.5 1691.1447692692693u,0 1693.0988493493492u,0 1693.0998493493494u,1.5 1695.0539294294292u,1.5 1695.0549294294294u,0 1696.0314694694694u,0 1696.0324694694696u,1.5 1698.9640895895895u,1.5 1698.9650895895898u,0 1701.8967097097095u,0 1701.8977097097097u,1.5 1702.8742497497497u,1.5 1702.8752497497499u,0 1705.8068698698698u,0 1705.80786986987u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1712.6496501501501u,0 1712.6506501501503u,1.5 1713.6271901901903u,1.5 1713.6281901901905u,0 1714.6047302302302u,0 1714.6057302302304u,1.5 1719.4924304304302u,1.5 1719.4934304304304u,0 1720.4699704704703u,0 1720.4709704704705u,1.5 1721.4475105105103u,1.5 1721.4485105105105u,0 1723.4025905905905u,0 1723.4035905905907u,1.5 1727.3127507507506u,1.5 1727.3137507507508u,0 1729.2678308308307u,0 1729.268830830831u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1735.133071071071u,0 1735.1340710710713u,1.5 1737.0881511511511u,1.5 1737.0891511511513u,0 1738.0656911911913u,0 1738.0666911911915u,1.5 1740.998311311311u,1.5 1740.9993113113112u,0 1741.9758513513511u,0 1741.9768513513513u,1.5 1742.9533913913913u,1.5 1742.9543913913915u,0 1745.8860115115112u,0 1745.8870115115114u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1754.6838718718718u,1.5 1754.684871871872u,0 1755.6614119119117u,0 1755.662411911912u,1.5 1758.594032032032u,1.5 1758.5950320320321u,0 1759.571572072072u,0 1759.5725720720723u,1.5 1761.526652152152u,1.5 1761.5276521521523u,0 1764.4592722722723u,0 1764.4602722722725u,1.5 1766.4143523523521u,1.5 1766.4153523523523u,0 1768.3694324324322u,0 1768.3704324324324u,1.5 1771.3020525525524u,1.5 1771.3030525525526u,0 1774.2346726726726u,0 1774.2356726726728u,1.5 1775.2122127127125u,1.5 1775.2132127127127u,0 1777.1672927927928u,0 1777.168292792793u,1.5 1779.1223728728728u,1.5 1779.123372872873u,0 1780.0999129129127u,0 1780.100912912913u,1.5 1781.0774529529529u,1.5 1781.078452952953u,0 1784.010073073073u,0 1784.0110730730732u,1.5 1784.987613113113u,1.5 1784.9886131131132u,0 1788.8977732732733u,0 1788.8987732732735u,1.5 1790.852853353353u,1.5 1790.8538533533533u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1794.7630135135132u,0 1794.7640135135134u,1.5 1796.7180935935935u,1.5 1796.7190935935937u,0 1798.6731736736735u,0 1798.6741736736737u,1.5 1802.5833338338336u,1.5 1802.5843338338339u,0 1803.5608738738738u,0 1803.561873873874u,1.5 1804.5384139139137u,1.5 1804.539413913914u,0 1807.471034034034u,0 1807.472034034034u,1.5 1808.448574074074u,1.5 1808.4495740740742u,0 1809.426114114114u,0 1809.4271141141141u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1820.1790545545543u,0 1820.1800545545545u,1.5 1821.1565945945945u,1.5 1821.1575945945947u,0 1822.1341346346344u,0 1822.1351346346346u,1.5 1823.1116746746745u,1.5 1823.1126746746747u,0 1824.0892147147147u,0 1824.0902147147149u,1.5 1826.0442947947947u,1.5 1826.045294794795u,0 1832.887075075075u,0 1832.8880750750752u,1.5 1834.842155155155u,1.5 1834.8431551551553u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1839.7298553553553u,1.5 1839.7308553553555u,0 1843.6400155155154u,0 1843.6410155155156u,1.5 1845.5950955955955u,1.5 1845.5960955955957u,0 1846.5726356356354u,0 1846.5736356356356u,1.5 1851.4603358358356u,1.5 1851.4613358358358u,0 1854.3929559559558u,0 1854.393955955956u,1.5 1857.325576076076u,1.5 1857.3265760760762u,0 1858.3031161161161u,0 1858.3041161161163u,1.5 1863.1908163163164u,1.5 1863.1918163163166u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1866.1234364364361u,1.5 1866.1244364364363u,0 1871.0111366366364u,0 1871.0121366366366u,1.5 1871.9886766766765u,1.5 1871.9896766766767u,0 1872.9662167167166u,0 1872.9672167167168u,1.5 1876.8763768768767u,1.5 1876.877376876877u,0 1877.853916916917u,0 1877.854916916917u,1.5 1878.8314569569568u,1.5 1878.832456956957u,0 1883.719157157157u,0 1883.7201571571572u,1.5 1884.6966971971972u,1.5 1884.6976971971974u,0 1885.674237237237u,0 1885.6752372372373u,1.5 1887.6293173173174u,1.5 1887.6303173173176u,0 1888.6068573573573u,0 1888.6078573573575u,1.5 1889.5843973973974u,1.5 1889.5853973973976u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1900.3373378378376u,1.5 1900.3383378378378u,0 1903.2699579579578u,0 1903.270957957958u,1.5 1905.2250380380378u,1.5 1905.226038038038u,0 1906.202578078078u,0 1906.2035780780782u,1.5 1908.157658158158u,1.5 1908.1586581581582u,0 1909.1351981981982u,0 1909.1361981981984u,1.5 1911.0902782782782u,1.5 1911.0912782782784u,0 1915.0004384384383u,0 1915.0014384384385u,1.5 1916.9555185185184u,1.5 1916.9565185185186u,0 1919.8881386386383u,0 1919.8891386386385u,1.5 1920.8656786786785u,1.5 1920.8666786786787u,0 1922.8207587587585u,0 1922.8217587587587u,1.5 1924.7758388388386u,1.5 1924.7768388388388u,0 1925.7533788788787u,0 1925.754378878879u,1.5 1926.7309189189189u,1.5 1926.731918918919u,0 1927.7084589589588u,0 1927.709458958959u,1.5 1929.6635390390388u,1.5 1929.664539039039u,0 1930.641079079079u,0 1930.6420790790792u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1940.4164794794794u,0 1940.4174794794797u,1.5 1942.3715595595593u,1.5 1942.3725595595595u,0 1943.3490995995994u,0 1943.3500995995996u,1.5 1946.2817197197196u,1.5 1946.2827197197198u,0 1948.2367997997997u,0 1948.2377997997999u,1.5 1949.2143398398398u,1.5 1949.21533983984u,0 1950.1918798798797u,0 1950.19287987988u,1.5 1951.1694199199198u,1.5 1951.17041991992u,0 1953.1245u,0 1953.1255u,1.5 1956.0571201201199u,1.5 1956.05812012012u,0 1957.03466016016u,0 1957.0356601601602u,1.5 1958.9897402402403u,1.5 1958.9907402402405u,0 1961.9223603603602u,0 1961.9233603603604u,1.5 1964.8549804804804u,1.5 1964.8559804804806u,0 1965.8325205205203u,0 1965.8335205205206u,1.5 1967.7876006006004u,1.5 1967.7886006006006u,0 1968.7651406406405u,0 1968.7661406406407u,1.5 1970.7202207207204u,1.5 1970.7212207207206u,0 1971.6977607607605u,0 1971.6987607607607u,1.5 1974.630380880881u,1.5 1974.6313808808811u,0 1976.5854609609607u,0 1976.586460960961u,1.5 1977.5630010010009u,1.5 1977.564001001001u,0 1980.4956211211208u,0 1980.496621121121u,1.5 1981.473161161161u,1.5 1981.4741611611612u,0 1983.4282412412413u,0 1983.4292412412415u,1.5 1984.4057812812814u,1.5 1984.4067812812816u,0 1986.3608613613612u,0 1986.3618613613614u,1.5 1991.2485615615612u,1.5 1991.2495615615614u,0 1992.2261016016014u,0 1992.2271016016016u,1.5 1993.2036416416415u,1.5 1993.2046416416417u,0 1995.1587217217213u,0 1995.1597217217216u,1.5 1997.1138018018016u,1.5 1997.1148018018018u,0 1998.0913418418418u,0 1998.092341841842u,1.5 1999.068881881882u,1.5 1999.069881881882u,0 2005.911662162162u,0 2005.9126621621622u,1.5 2006.8892022022021u,1.5 2006.8902022022023u,0 2007.8667422422423u,0 2007.8677422422425u,1.5 2009.821822322322u,1.5 2009.8228223223223u,0 2014.7095225225223u,0 2014.7105225225225u,1.5 2015.6870625625625u,1.5 2015.6880625625627u,0 2021.5523028028026u,0 2021.5533028028028u,1.5 2022.5298428428428u,1.5 2022.530842842843u,0 2023.507382882883u,0 2023.508382882883u,1.5 2024.4849229229226u,1.5 2024.4859229229228u,0 2025.4624629629627u,0 2025.463462962963u,1.5 2026.4400030030029u,1.5 2026.441003003003u,0 2027.417543043043u,0 2027.4185430430432u,1.5 2028.3950830830831u,1.5 2028.3960830830833u,0 2029.3726231231228u,0 2029.373623123123u,1.5 2032.3052432432432u,1.5 2032.3062432432434u,0 2033.2827832832834u,0 2033.2837832832836u,1.5 2036.2154034034033u,1.5 2036.2164034034035u,0 2037.1929434434435u,0 2037.1939434434437u,1.5 2040.1255635635634u,1.5 2040.1265635635636u,0 2042.0806436436435u,0 2042.0816436436437u,1.5 2043.0581836836836u,1.5 2043.0591836836838u,0 2044.0357237237233u,0 2044.0367237237235u,1.5 2046.9683438438437u,1.5 2046.969343843844u,0 2047.9458838838839u,0 2047.946883883884u,1.5 2048.9234239239236u,1.5 2048.9244239239238u,0 2049.900963963964u,0 2049.901963963964u,1.5 2051.856044044044u,1.5 2051.8570440440444u,0 2054.788664164164u,0 2054.789664164164u,1.5 2055.766204204204u,1.5 2055.767204204204u,0 2058.698824324324u,0 2058.6998243243243u,1.5 2060.6539044044043u,1.5 2060.6549044044045u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2067.4966846846846u,0 2067.497684684685u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2070.429304804805u,0 2070.430304804805u,1.5 2074.339464964965u,1.5 2074.340464964965u,0 2075.317005005005u,0 2075.318005005005u,1.5 2077.272085085085u,1.5 2077.2730850850853u,0 2078.249625125125u,0 2078.250625125125u,1.5 2079.227165165165u,1.5 2079.228165165165u,0 2086.0699454454452u,0 2086.0709454454454u,1.5 2091.9351856856856u,1.5 2091.936185685686u,0 2092.9127257257255u,0 2092.9137257257257u,1.5 2095.8453458458457u,1.5 2095.846345845846u,0 2096.822885885886u,0 2096.8238858858863u,1.5 2097.8004259259255u,1.5 2097.8014259259257u,0 2102.688126126126u,0 2102.689126126126u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2105.620746246246u,0 2105.6217462462464u,1.5 2114.4186066066063u,1.5 2114.4196066066065u,0 2120.2838468468467u,0 2120.284846846847u,1.5 2121.261386886887u,1.5 2121.2623868868873u,0 2123.216466966967u,0 2123.217466966967u,1.5 2127.126627127127u,1.5 2127.127627127127u,0 2128.104167167167u,0 2128.105167167167u,1.5 2129.081707207207u,1.5 2129.082707207207u,0 2132.991867367367u,0 2132.992867367367u,1.5 2133.9694074074073u,1.5 2133.9704074074075u,0 2134.946947447447u,0 2134.9479474474474u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2137.8795675675674u,0 2137.8805675675676u,1.5 2138.8571076076073u,1.5 2138.8581076076075u,0 2140.8121876876876u,0 2140.813187687688u,1.5 2142.7672677677674u,1.5 2142.7682677677676u,0 2143.744807807808u,0 2143.745807807808u,1.5 2144.7223478478477u,1.5 2144.723347847848u,0 2145.699887887888u,0 2145.7008878878883u,1.5 2146.677427927928u,1.5 2146.678427927928u,0 2149.610048048048u,0 2149.6110480480484u,1.5 2154.497748248248u,1.5 2154.4987482482484u,0 2156.4528283283285u,0 2156.4538283283287u,1.5 2157.430368368368u,1.5 2157.431368368368u,0 2162.3180685685684u,0 2162.3190685685686u,1.5 2163.2956086086083u,1.5 2163.2966086086085u,0 2164.2731486486487u,0 2164.274148648649u,1.5 2167.2057687687684u,1.5 2167.2067687687686u,0 2169.1608488488487u,0 2169.161848848849u,1.5 2170.138388888889u,1.5 2170.1393888888892u,0 2174.048549049049u,0 2174.0495490490493u,1.5 2180.8913293293294u,1.5 2180.8923293293296u,0 2181.868869369369u,0 2181.869869369369u,1.5 2182.8464094094093u,1.5 2182.8474094094095u,0 2184.8014894894895u,0 2184.8024894894897u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2187.7341096096093u,0 2187.7351096096095u,1.5 2191.6442697697694u,1.5 2191.6452697697696u,0 2196.53196996997u,0 2196.53296996997u,1.5 2197.5095100100098u,1.5 2197.51051001001u,0 2198.48705005005u,0 2198.4880500500503u,1.5 2200.4421301301304u,1.5 2200.4431301301306u,0 2201.41967017017u,0 2201.42067017017u,1.5 2203.37475025025u,1.5 2203.3757502502503u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2211.1950705705704u,1.5 2211.1960705705706u,0 2212.1726106106103u,0 2212.1736106106105u,1.5 2215.105230730731u,1.5 2215.106230730731u,0 2219.992930930931u,0 2219.993930930931u,1.5 2220.970470970971u,1.5 2220.971470970971u,0 2221.9480110110107u,0 2221.949011011011u,1.5 2223.903091091091u,1.5 2223.9040910910912u,0 2227.813251251251u,0 2227.8142512512513u,1.5 2228.790791291291u,1.5 2228.7917912912912u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2230.745871371371u,1.5 2230.746871371371u,0 2232.700951451451u,0 2232.7019514514514u,1.5 2234.6560315315314u,1.5 2234.6570315315316u,0 2235.6335715715713u,0 2235.6345715715715u,1.5 2236.6111116116112u,1.5 2236.6121116116115u,0 2238.5661916916915u,0 2238.5671916916917u,1.5 2239.543731731732u,1.5 2239.544731731732u,0 2240.5212717717714u,0 2240.5222717717716u,1.5 2241.4988118118117u,1.5 2241.499811811812u,0 2242.4763518518516u,0 2242.477351851852u,1.5 2243.453891891892u,1.5 2243.454891891892u,0 2244.431431931932u,0 2244.432431931932u,1.5 2245.408971971972u,1.5 2245.409971971972u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2255.184372372372u,0 2255.185372372372u,1.5 2256.161912412412u,1.5 2256.1629124124124u,0 2260.0720725725723u,0 2260.0730725725725u,1.5 2264.9597727727723u,1.5 2264.9607727727725u,0 2265.9373128128127u,0 2265.938312812813u,1.5 2266.9148528528526u,1.5 2266.915852852853u,0 2267.892392892893u,0 2267.893392892893u,1.5 2269.847472972973u,1.5 2269.848472972973u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2276.690253253253u,1.5 2276.6912532532533u,0 2277.6677932932935u,0 2277.6687932932937u,1.5 2278.6453333333334u,1.5 2278.6463333333336u,0 2280.600413413413u,0 2280.6014134134134u,1.5 2281.577953453453u,1.5 2281.5789534534533u,0 2282.5554934934935u,0 2282.5564934934937u,1.5 2284.5105735735733u,1.5 2284.5115735735735u,0 2285.488113613613u,0 2285.4891136136134u,1.5 2287.4431936936935u,1.5 2287.4441936936937u,0 2288.420733733734u,0 2288.421733733734u,1.5 2289.3982737737733u,1.5 2289.3992737737735u,0 2290.3758138138137u,0 2290.376813813814u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2293.308433933934u,0 2293.309433933934u,1.5 2299.173674174174u,1.5 2299.174674174174u,0 2304.0613743743743u,0 2304.0623743743745u,1.5 2307.9715345345344u,1.5 2307.9725345345346u,0 2308.9490745745743u,0 2308.9500745745745u,1.5 2309.926614614614u,1.5 2309.9276146146144u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2314.8143148148147u,1.5 2314.815314814815u,0 2319.7020150150147u,0 2319.703015015015u,1.5 2320.679555055055u,1.5 2320.6805550550553u,0 2324.589715215215u,0 2324.5907152152154u,1.5 2325.567255255255u,1.5 2325.5682552552553u,0 2327.5223353353354u,0 2327.5233353353356u,1.5 2332.4100355355354u,1.5 2332.4110355355356u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2340.2303558558556u,1.5 2340.231355855856u,0 2341.207895895896u,0 2341.208895895896u,1.5 2342.185435935936u,1.5 2342.186435935936u,0 2343.1629759759758u,0 2343.163975975976u,1.5 2344.1405160160157u,1.5 2344.141516016016u,0 2349.028216216216u,0 2349.0292162162164u,1.5 2350.005756256256u,1.5 2350.0067562562563u,0 2350.9832962962964u,0 2350.9842962962966u,1.5 2354.893456456456u,1.5 2354.8944564564563u,0 2355.8709964964964u,0 2355.8719964964966u,1.5 2356.8485365365364u,1.5 2356.8495365365366u,0 2358.803616616616u,0 2358.8046166166164u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2366.623936936937u,0 2366.624936936937u,1.5 2367.6014769769768u,1.5 2367.602476976977u,0 2369.556557057057u,0 2369.5575570570572u,1.5 2371.5116371371373u,1.5 2371.5126371371375u,0 2376.3993373373373u,0 2376.4003373373375u,1.5 2377.3768773773777u,1.5 2377.377877377378u,0 2380.3094974974974u,0 2380.3104974974976u,1.5 2386.174737737738u,1.5 2386.175737737738u,0 2387.1522777777777u,0 2387.153277777778u,1.5 2388.1298178178176u,1.5 2388.130817817818u,0 2393.995058058058u,0 2393.996058058058u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2398.882758258258u,0 2398.8837582582582u,1.5 2400.8378383383383u,1.5 2400.8388383383385u,0 2401.8153783783787u,0 2401.816378378379u,1.5 2402.792918418418u,1.5 2402.7939184184183u,0 2403.7704584584585u,0 2403.7714584584587u,1.5 2405.7255385385383u,1.5 2405.7265385385385u,0 2410.613238738739u,0 2410.614238738739u,1.5 2411.5907787787787u,1.5 2411.591778778779u,0 2412.5683188188186u,0 2412.569318818819u,1.5 2415.500938938939u,1.5 2415.501938938939u,0 2416.478478978979u,0 2416.4794789789794u,1.5 2423.321259259259u,1.5 2423.322259259259u,0 2425.2763393393393u,0 2425.2773393393395u,1.5 2426.2538793793797u,1.5 2426.25487937938u,0 2432.119119619619u,0 2432.1201196196193u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2435.05173973974u,1.5 2435.05273973974u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.9843598598595u,1.5 2437.9853598598597u,0 2438.9618998999u,0 2438.9628998999u,1.5 2441.8945200200196u,1.5 2441.89552002002u,0 2442.87206006006u,0 2442.87306006006u,1.5 2446.78222022022u,1.5 2446.7832202202203u,0 2447.75976026026u,0 2447.76076026026u,1.5 2449.7148403403403u,1.5 2449.7158403403405u,0 2451.66992042042u,0 2451.6709204204203u,1.5 2452.6474604604605u,1.5 2452.6484604604607u,0 2454.6025405405403u,0 2454.6035405405405u,1.5 2455.5800805805807u,1.5 2455.581080580581u,0 2459.490240740741u,0 2459.491240740741u,1.5 2462.4228608608605u,1.5 2462.4238608608607u,0 2464.377940940941u,0 2464.378940940941u,1.5 2465.355480980981u,1.5 2465.3564809809814u,0 2466.3330210210206u,0 2466.334021021021u,1.5 2467.310561061061u,1.5 2467.311561061061u,0 2468.288101101101u,0 2468.289101101101u,1.5 2472.198261261261u,1.5 2472.199261261261u,0 2474.1533413413413u,0 2474.1543413413415u,1.5 2476.108421421421u,1.5 2476.1094214214213u,0 2478.0635015015014u,0 2478.0645015015016u,1.5 2482.9512017017014u,1.5 2482.9522017017016u,0 2483.9287417417418u,0 2483.929741741742u,1.5 2484.9062817817817u,1.5 2484.907281781782u,0 2485.8838218218216u,0 2485.884821821822u,1.5 2500.546922422422u,1.5 2500.5479224224223u,0 2505.434622622622u,0 2505.4356226226223u,1.5 2512.277402902903u,1.5 2512.278402902903u,0 2513.2549429429428u,0 2513.255942942943u,1.5 2517.165103103103u,1.5 2517.166103103103u,0 2518.1426431431432u,0 2518.1436431431434u,1.5 2519.120183183183u,1.5 2519.1211831831833u,0 2520.097723223223u,0 2520.0987232232233u,1.5 2522.0528033033033u,1.5 2522.0538033033035u,0 2523.0303433433432u,0 2523.0313433433435u,1.5 2524.985423423423u,1.5 2524.9864234234233u,0 2525.9629634634634u,0 2525.9639634634636u,1.5 2527.9180435435437u,1.5 2527.919043543544u,0 2528.8955835835836u,0 2528.896583583584u,1.5 2529.8731236236235u,1.5 2529.8741236236237u,0 2531.8282037037034u,0 2531.8292037037036u,1.5 2532.8057437437437u,1.5 2532.806743743744u,0 2533.7832837837836u,0 2533.784283783784u,1.5 2534.7608238238236u,1.5 2534.7618238238238u,0 2539.6485240240236u,0 2539.649524024024u,1.5 2540.626064064064u,1.5 2540.627064064064u,0 2544.536224224224u,0 2544.5372242242242u,1.5 2546.4913043043043u,1.5 2546.4923043043045u,0 2547.4688443443442u,0 2547.4698443443444u,1.5 2548.4463843843846u,1.5 2548.447384384385u,0 2549.423924424424u,0 2549.4249244244243u,1.5 2550.4014644644644u,1.5 2550.4024644644646u,0 2552.3565445445447u,0 2552.357544544545u,1.5 2554.3116246246245u,1.5 2554.3126246246247u,0 2556.2667047047044u,0 2556.2677047047046u,1.5 2557.2442447447447u,1.5 2557.245244744745u,0 2562.1319449449447u,0 2562.132944944945u,1.5 2565.064565065065u,1.5 2565.065565065065u,0 2566.042105105105u,0 2566.043105105105u,1.5 2567.019645145145u,1.5 2567.0206451451454u,0 2567.997185185185u,0 2567.9981851851853u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2577.7725855855856u,0 2577.773585585586u,1.5 2586.5704459459457u,1.5 2586.571445945946u,0 2587.547985985986u,0 2587.5489859859863u,1.5 2588.5255260260255u,1.5 2588.5265260260257u,0 2596.345846346346u,0 2596.3468463463464u,1.5 2597.3233863863866u,1.5 2597.324386386387u,0 2598.300926426426u,0 2598.3019264264262u,1.5 2599.2784664664664u,1.5 2599.2794664664666u,0 2600.2560065065063u,0 2600.2570065065065u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2608.0763268268265u,1.5 2608.0773268268267u,0 2611.0089469469467u,0 2611.009946946947u,1.5 2611.986486986987u,1.5 2611.9874869869873u,0 2612.9640270270265u,0 2612.9650270270267u,1.5 2613.941567067067u,1.5 2613.942567067067u,0 2615.896647147147u,0 2615.8976471471474u,1.5 2619.8068073073073u,1.5 2619.8078073073075u,0 2620.784347347347u,0 2620.7853473473474u,1.5 2622.739427427427u,1.5 2622.740427427427u,0 2628.6046676676674u,0 2628.6056676676676u,1.5 2629.5822077077073u,1.5 2629.5832077077075u,0 2630.5597477477477u,0 2630.560747747748u,1.5 2634.469907907908u,1.5 2634.470907907908u,0 2635.4474479479477u,0 2635.448447947948u,1.5 2637.402528028028u,1.5 2637.403528028028u,0 2642.2902282282284u,0 2642.2912282282286u,1.5 2643.267768268268u,1.5 2643.268768268268u,0 2644.2453083083083u,0 2644.2463083083085u,1.5 2651.0880885885886u,1.5 2651.0890885885888u,0 2652.065628628629u,0 2652.066628628629u,1.5 2653.0431686686684u,1.5 2653.0441686686686u,0 2654.9982487487487u,0 2654.999248748749u,1.5 2655.9757887887886u,1.5 2655.976788788789u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2666.7287292292294u,1.5 2666.7297292292296u,0 2667.706269269269u,0 2667.707269269269u,1.5 2672.5939694694694u,1.5 2672.5949694694696u,0 2673.5715095095093u,0 2673.5725095095095u,1.5 2674.5490495495496u,1.5 2674.55004954955u,0 2679.4367497497497u,0 2679.43774974975u,1.5 2681.39182982983u,1.5 2681.39282982983u,0 2682.3693698698694u,0 2682.3703698698696u,1.5 2684.3244499499497u,1.5 2684.32544994995u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2689.21215015015u,0 2689.2131501501503u,1.5 2691.1672302302304u,1.5 2691.1682302302306u,0 2693.1223103103102u,0 2693.1233103103104u,1.5 2694.09985035035u,1.5 2694.1008503503504u,0 2695.0773903903905u,0 2695.0783903903907u,1.5 2696.0549304304304u,1.5 2696.0559304304306u,0 2698.0100105105103u,0 2698.0110105105105u,1.5 2698.9875505505506u,1.5 2698.988550550551u,0 2699.9650905905905u,0 2699.9660905905907u,1.5 2701.9201706706704u,1.5 2701.9211706706706u,0 2703.8752507507506u,0 2703.876250750751u,1.5 2706.8078708708704u,1.5 2706.8088708708706u,0 2710.718031031031u,0 2710.719031031031u,1.5 2713.650651151151u,1.5 2713.6516511511513u,0 2714.628191191191u,0 2714.6291911911912u,1.5 2718.538351351351u,1.5 2718.5393513513513u,0 2719.5158913913915u,0 2719.5168913913917u,1.5 2721.4709714714713u,1.5 2721.4719714714715u,0 2722.4485115115112u,0 2722.4495115115114u,1.5 2723.4260515515516u,1.5 2723.427051551552u,0 2725.381131631632u,0 2725.382131631632u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2730.268831831832u,1.5 2730.269831831832u,0 2733.2014519519516u,0 2733.202451951952u,1.5 2735.156532032032u,1.5 2735.157532032032u,0 2736.134072072072u,0 2736.135072072072u,1.5 2737.1116121121117u,1.5 2737.112612112112u,0 2738.089152152152u,0 2738.0901521521523u,1.5 2739.066692192192u,1.5 2739.067692192192u,0 2740.0442322322324u,0 2740.0452322322326u,1.5 2741.021772272272u,1.5 2741.022772272272u,0 2745.9094724724723u,0 2745.9104724724725u,1.5 2746.8870125125122u,1.5 2746.8880125125124u,0 2747.8645525525526u,0 2747.865552552553u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 2755.6848728728723u,0 2755.6858728728726u,1.5 2756.6624129129127u,1.5 2756.663412912913u,0 2757.6399529529526u,0 2757.640952952953u,1.5 2760.572573073073u,1.5 2760.573573073073u,0 2761.5501131131127u,0 2761.551113113113u,1.5 2762.527653153153u,1.5 2762.5286531531533u,0 2765.460273273273u,0 2765.461273273273u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2773.2805935935935u,1.5 2773.2815935935937u,0 2777.1907537537536u,0 2777.191753753754u,1.5 2782.0784539539536u,1.5 2782.079453953954u,0 2786.966154154154u,0 2786.9671541541543u,1.5 2787.943694194194u,1.5 2787.944694194194u,0 2788.9212342342344u,0 2788.9222342342346u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2795.764014514514u,0 2795.7650145145144u,1.5 2796.7415545545546u,1.5 2796.7425545545548u,0 2798.696634634635u,0 2798.697634634635u,1.5 2800.6517147147147u,1.5 2800.652714714715u,0 2803.584334834835u,0 2803.585334834835u,1.5 2804.561874874875u,1.5 2804.562874874875u,0 2805.5394149149147u,0 2805.540414914915u,1.5 2806.5169549549546u,1.5 2806.517954954955u,0 2808.472035035035u,0 2808.473035035035u,1.5 2809.449575075075u,1.5 2809.450575075075u,0 2810.4271151151147u,0 2810.428115115115u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2819.2249754754753u,0 2819.2259754754755u,1.5 2820.202515515515u,1.5 2820.2035155155154u,0 2829.9779159159157u,0 2829.978915915916u,1.5 2831.932995995996u,1.5 2831.933995995996u,0 2833.888076076076u,0 2833.889076076076u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2839.753316316316u,0 2839.7543163163164u,1.5 2840.730856356356u,1.5 2840.7318563563563u,0 2844.641016516516u,0 2844.6420165165164u,1.5 2846.5960965965965u,1.5 2846.5970965965967u,0 2847.573636636637u,0 2847.574636636637u,1.5 2848.5511766766763u,1.5 2848.5521766766765u,0 2850.5062567567566u,0 2850.5072567567568u,1.5 2852.461336836837u,1.5 2852.462336836837u,0 2855.3939569569566u,0 2855.394956956957u,1.5 2856.371496996997u,1.5 2856.372496996997u,0 2857.349037037037u,0 2857.350037037037u,1.5 2859.3041171171167u,1.5 2859.305117117117u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2865.169357357357u,0 2865.1703573573573u,1.5 2866.1468973973974u,1.5 2866.1478973973976u,0 2871.0345975975974u,0 2871.0355975975976u,1.5 2874.9447577577575u,1.5 2874.9457577577577u,0 2876.899837837838u,0 2876.900837837838u,1.5 2877.877377877878u,1.5 2877.8783778778784u,0 2878.8549179179176u,0 2878.855917917918u,1.5 2879.832457957958u,1.5 2879.833457957958u,0 2880.809997997998u,0 2880.810997997998u,1.5 2881.787538038038u,1.5 2881.788538038038u,0 2882.765078078078u,0 2882.7660780780784u,1.5 2883.7426181181177u,1.5 2883.743618118118u,0 2885.697698198198u,0 2885.698698198198u,1.5 2886.6752382382383u,1.5 2886.6762382382385u,0 2887.652778278278u,0 2887.6537782782784u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2899.3832587587585u,0 2899.3842587587587u,1.5 2900.360798798799u,1.5 2900.361798798799u,0 2901.338338838839u,0 2901.339338838839u,1.5 2902.315878878879u,1.5 2902.3168788788794u,0 2903.2934189189186u,0 2903.294418918919u,1.5 2909.158659159159u,1.5 2909.159659159159u,0 2910.136199199199u,0 2910.137199199199u,1.5 2912.091279279279u,1.5 2912.0922792792794u,0 2913.068819319319u,0 2913.0698193193193u,1.5 2914.046359359359u,1.5 2914.0473593593592u,0 2921.8666796796797u,0 2921.86767967968u,1.5 2922.8442197197196u,1.5 2922.84521971972u,0 2923.8217597597595u,0 2923.8227597597597u,1.5 2930.66454004004u,1.5 2930.66554004004u,0 2931.64208008008u,0 2931.6430800800804u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2938.48486036036u,0 2938.48586036036u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 2946.3051806806807u,0 2946.306180680681u,1.5 2947.2827207207206u,1.5 2947.283720720721u,0 2948.2602607607605u,0 2948.2612607607607u,1.5 2949.237800800801u,1.5 2949.238800800801u,0 2950.215340840841u,0 2950.216340840841u,1.5 2955.103041041041u,1.5 2955.104041041041u,0 2956.080581081081u,0 2956.0815810810814u,1.5 2958.035661161161u,1.5 2958.036661161161u,0 2959.013201201201u,0 2959.014201201201u,1.5 2962.923361361361u,1.5 2962.924361361361u,0 2963.9009014014014u,0 2963.9019014014016u,1.5 2965.8559814814816u,1.5 2965.856981481482u,0 2966.833521521521u,0 2966.8345215215213u,1.5 2968.7886016016014u,1.5 2968.7896016016016u,0 2969.7661416416418u,0 2969.767141641642u,1.5 2970.7436816816817u,1.5 2970.744681681682u,0 2971.7212217217216u,0 2971.722221721722u,1.5 2972.6987617617615u,1.5 2972.6997617617617u,0 2973.676301801802u,0 2973.677301801802u,1.5 2974.6538418418418u,1.5 2974.654841841842u,0 2979.541542042042u,0 2979.542542042042u,1.5 2980.519082082082u,1.5 2980.5200820820824u,0 2982.474162162162u,0 2982.475162162162u,1.5 2983.451702202202u,1.5 2983.452702202202u,0 2992.2495625625625u,0 2992.2505625625627u,1.5 2993.2271026026024u,1.5 2993.2281026026026u,0 2999.0923428428428u,0 2999.093342842843u,1.5 3000.069882882883u,1.5 3000.0708828828833u,0 3003.002503003003u,0 3003.003503003003u,1.5 3003.980043043043u,1.5 3003.9810430430434u,0 3006.912663163163u,0 3006.913663163163u,1.5 3009.845283283283u,1.5 3009.8462832832834u,0 3010.822823323323u,0 3010.8238233233233u,1.5 3011.800363363363u,1.5 3011.801363363363u,0 3013.7554434434433u,0 3013.7564434434435u,1.5 3014.7329834834836u,1.5 3014.733983483484u,0 3016.6880635635634u,0 3016.6890635635636u,1.5 3017.6656036036034u,1.5 3017.6666036036036u,0 3018.6431436436437u,0 3018.644143643644u,1.5 3019.6206836836836u,1.5 3019.621683683684u,0 3022.553303803804u,0 3022.554303803804u,1.5 3024.508383883884u,1.5 3024.5093838838843u,0 3025.4859239239236u,0 3025.4869239239238u,1.5 3027.441004004004u,1.5 3027.442004004004u,0 3028.418544044044u,0 3028.4195440440444u,1.5 3029.396084084084u,1.5 3029.3970840840843u,0 3030.373624124124u,0 3030.3746241241242u,1.5 3032.328704204204u,1.5 3032.329704204204u,0 3033.306244244244u,0 3033.3072442442444u,1.5 3034.283784284284u,1.5 3034.2847842842843u,0 3035.261324324324u,0 3035.2623243243243u,1.5 3038.1939444444442u,1.5 3038.1949444444444u,0 3039.1714844844846u,0 3039.172484484485u,1.5 3040.149024524524u,1.5 3040.1500245245243u,0 3041.1265645645644u,0 3041.1275645645646u,1.5 3042.1041046046043u,1.5 3042.1051046046045u,0 3044.0591846846846u,0 3044.060184684685u,1.5 3046.0142647647644u,1.5 3046.0152647647647u,0 3046.991804804805u,0 3046.992804804805u,1.5 3048.946884884885u,1.5 3048.9478848848853u,0 3050.901964964965u,0 3050.902964964965u,1.5 3052.857045045045u,1.5 3052.8580450450454u,0 3054.812125125125u,0 3054.813125125125u,1.5 3055.789665165165u,1.5 3055.790665165165u,0 3062.6324454454452u,0 3062.6334454454454u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3066.5426056056053u,1.5 3066.5436056056055u,0 3067.5201456456457u,0 3067.521145645646u,1.5 3073.385385885886u,1.5 3073.3863858858863u,0 3074.3629259259255u,0 3074.3639259259257u,1.5 3077.295546046046u,1.5 3077.2965460460464u,0 3079.250626126126u,0 3079.251626126126u,1.5 3080.228166166166u,1.5 3080.229166166166u,0 3084.138326326326u,0 3084.139326326326u,1.5 3085.115866366366u,1.5 3085.116866366366u,0 3088.0484864864866u,0 3088.049486486487u,1.5 3090.0035665665664u,1.5 3090.0045665665666u,0 3090.9811066066063u,0 3090.9821066066065u,1.5 3092.9361866866866u,1.5 3092.937186686687u,0 3093.9137267267265u,0 3093.9147267267267u,1.5 3094.8912667667664u,1.5 3094.8922667667666u,0 3095.868806806807u,0 3095.869806806807u,1.5 3096.8463468468467u,1.5 3096.847346846847u,0 3097.823886886887u,0 3097.8248868868873u,1.5 3098.8014269269265u,1.5 3098.8024269269267u,0 3102.711587087087u,0 3102.7125870870873u,1.5 3104.666667167167u,1.5 3104.667667167167u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3112.4869874874876u,1.5 3112.4879874874878u,0 3113.464527527527u,0 3113.4655275275272u,1.5 3114.4420675675674u,1.5 3114.4430675675676u,0 3115.4196076076073u,0 3115.4206076076075u,1.5 3116.3971476476477u,1.5 3116.398147647648u,0 3118.3522277277275u,0 3118.3532277277277u,1.5 3120.307307807808u,1.5 3120.308307807808u,0 3122.262387887888u,0 3122.2633878878883u,1.5 3125.195008008008u,1.5 3125.196008008008u,0 3126.172548048048u,0 3126.1735480480484u,1.5 3127.150088088088u,1.5 3127.1510880880883u,0 3128.127628128128u,0 3128.128628128128u,1.5 3131.060248248248u,1.5 3131.0612482482484u,0 3135.947948448448u,0 3135.9489484484484u,1.5 3139.8581086086083u,1.5 3139.8591086086085u,0 3140.8356486486487u,0 3140.836648648649u,1.5 3143.7682687687684u,1.5 3143.7692687687686u,0 3147.678428928929u,0 3147.679428928929u,1.5 3148.655968968969u,1.5 3148.656968968969u,0 3151.588589089089u,0 3151.5895890890893u,1.5 3153.543669169169u,1.5 3153.544669169169u,0 3154.5212092092092u,0 3154.5222092092094u,1.5 3155.498749249249u,1.5 3155.4997492492494u,0 3156.476289289289u,0 3156.4772892892893u,1.5 3157.4538293293294u,1.5 3157.4548293293296u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3168.2067697697694u,1.5 3168.2077697697696u,0 3169.1843098098097u,0 3169.18530980981u,1.5 3170.1618498498497u,1.5 3170.16284984985u,0 3175.04955005005u,0 3175.0505500500503u,1.5 3177.0046301301304u,1.5 3177.0056301301306u,0 3178.9597102102102u,0 3178.9607102102104u,1.5 3179.93725025025u,1.5 3179.9382502502503u,0 3180.91479029029u,0 3180.9157902902903u,1.5 3182.86987037037u,1.5 3182.87087037037u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3190.6901906906905u,1.5 3190.6911906906907u,0 3191.667730730731u,0 3191.668730730731u,1.5 3192.6452707707704u,1.5 3192.6462707707706u,0 3196.555430930931u,0 3196.556430930931u,1.5 3197.532970970971u,1.5 3197.533970970971u,0 3198.5105110110107u,0 3198.511511011011u,1.5 3202.420671171171u,1.5 3202.421671171171u,0 3203.398211211211u,0 3203.3992112112114u,1.5 3204.375751251251u,1.5 3204.3767512512513u,0 3207.308371371371u,0 3207.309371371371u,1.5 3213.1736116116112u,1.5 3213.1746116116115u,0 3215.1286916916915u,0 3215.1296916916917u,1.5 3217.0837717717714u,1.5 3217.0847717717716u,0 3218.0613118118117u,0 3218.062311811812u,1.5 3219.0388518518516u,1.5 3219.039851851852u,0 3220.016391891892u,0 3220.017391891892u,1.5 3223.926552052052u,1.5 3223.9275520520523u,0 3224.904092092092u,0 3224.905092092092u,1.5 3225.8816321321324u,1.5 3225.8826321321326u,0 3227.836712212212u,0 3227.8377122122124u,1.5 3228.814252252252u,1.5 3228.8152522522523u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3232.724412412412u,1.5 3232.7254124124124u,0 3234.6794924924925u,0 3234.6804924924927u,1.5 3236.6345725725723u,1.5 3236.6355725725725u,0 3237.6121126126122u,0 3237.6131126126124u,1.5 3238.5896526526526u,1.5 3238.590652652653u,0 3239.5671926926925u,0 3239.5681926926927u,1.5 3240.544732732733u,1.5 3240.545732732733u,0 3242.4998128128127u,0 3242.500812812813u,1.5 3244.454892892893u,1.5 3244.455892892893u,0 3245.432432932933u,0 3245.433432932933u,1.5 3246.409972972973u,1.5 3246.410972972973u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3255.2078333333334u,1.5 3255.2088333333336u,0 3259.1179934934935u,0 3259.1189934934937u,1.5 3260.0955335335334u,1.5 3260.0965335335336u,0 3262.050613613613u,0 3262.0516136136134u,1.5 3263.0281536536536u,1.5 3263.029153653654u,0 3264.0056936936935u,0 3264.0066936936937u,1.5 3264.983233733734u,1.5 3264.984233733734u,0 3265.9607737737733u,0 3265.9617737737735u,1.5 3267.9158538538536u,1.5 3267.916853853854u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3274.7586341341344u,0 3274.7596341341346u,1.5 3277.691254254254u,1.5 3277.6922542542543u,0 3278.6687942942945u,0 3278.6697942942947u,1.5 3279.6463343343344u,1.5 3279.6473343343346u,0 3280.6238743743743u,0 3280.6248743743745u,1.5 3281.601414414414u,1.5 3281.6024144144144u,0 3283.5564944944945u,0 3283.5574944944947u,1.5 3285.5115745745743u,1.5 3285.5125745745745u,0 3286.489114614614u,0 3286.4901146146144u,1.5 3287.4666546546546u,1.5 3287.467654654655u,0 3289.421734734735u,0 3289.422734734735u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3294.309434934935u,0 3294.310434934935u,1.5 3297.242055055055u,1.5 3297.2430550550553u,0 3298.219595095095u,0 3298.220595095095u,1.5 3299.1971351351353u,1.5 3299.1981351351355u,0 3302.129755255255u,0 3302.1307552552553u,1.5 3303.1072952952954u,1.5 3303.1082952952956u,0 3304.0848353353354u,0 3304.0858353353356u,1.5 3307.9949954954955u,1.5 3307.9959954954957u,0 3308.9725355355354u,0 3308.9735355355356u,1.5 3310.927615615615u,1.5 3310.9286156156154u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3320.7030160160157u,1.5 3320.704016016016u,0 3325.590716216216u,0 3325.5917162162164u,1.5 3330.478416416416u,1.5 3330.4794164164164u,0 3331.455956456456u,0 3331.4569564564563u,1.5 3332.4334964964964u,1.5 3332.4344964964966u,0 3334.3885765765763u,0 3334.3895765765765u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3345.1415170170167u,1.5 3345.142517017017u,0 3347.096597097097u,0 3347.097597097097u,1.5 3348.0741371371373u,1.5 3348.0751371371375u,0 3349.0516771771768u,0 3349.052677177177u,1.5 3350.029217217217u,1.5 3350.0302172172173u,0 3351.006757257257u,0 3351.0077572572573u,1.5 3351.9842972972974u,1.5 3351.9852972972976u,0 3352.9618373373373u,0 3352.9628373373375u,1.5 3353.9393773773772u,1.5 3353.9403773773774u,0 3355.894457457457u,0 3355.8954574574573u,1.5 3357.8495375375373u,1.5 3357.8505375375375u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3365.6698578578576u,1.5 3365.6708578578578u,0 3366.647397897898u,0 3366.648397897898u,1.5 3369.5800180180177u,1.5 3369.581018018018u,0 3370.557558058058u,0 3370.558558058058u,1.5 3371.535098098098u,1.5 3371.536098098098u,0 3378.3778783783787u,0 3378.378878378379u,1.5 3382.2880385385383u,1.5 3382.2890385385385u,0 3384.243118618618u,0 3384.2441186186184u,1.5 3385.2206586586585u,1.5 3385.2216586586587u,0 3386.1981986986984u,0 3386.1991986986986u,1.5 3387.175738738739u,1.5 3387.176738738739u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3390.1083588588585u,1.5 3390.1093588588587u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3396.9511391391393u,0 3396.9521391391395u,1.5 3401.8388393393393u,1.5 3401.8398393393395u,0 3402.8163793793797u,0 3402.81737937938u,1.5 3404.7714594594595u,1.5 3404.7724594594597u,0 3409.6591596596595u,0 3409.6601596596597u,1.5 3410.6366996996994u,1.5 3410.6376996996996u,0 3413.5693198198196u,0 3413.57031981982u,1.5 3414.5468598598595u,1.5 3414.5478598598597u,0 3419.43456006006u,0 3419.43556006006u,1.5 3420.4121001001u,1.5 3420.4131001001u,0 3421.3896401401403u,0 3421.3906401401405u,1.5 3422.36718018018u,1.5 3422.3681801801804u,0 3423.34472022022u,0 3423.3457202202203u,1.5 3424.32226026026u,1.5 3424.32326026026u,0 3426.2773403403403u,0 3426.2783403403405u,1.5 3427.2548803803807u,1.5 3427.255880380381u,0 3430.1875005005004u,0 3430.1885005005006u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3434.0976606606605u,0 3434.0986606606607u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3436.052740740741u,0 3436.053740740741u,1.5 3450.7158413413413u,1.5 3450.7168413413415u,0 3451.6933813813816u,0 3451.694381381382u,1.5 3452.670921421421u,1.5 3452.6719214214213u,0 3454.6260015015014u,0 3454.6270015015016u,1.5 3457.558621621621u,1.5 3457.5596216216213u,0 3458.5361616616615u,0 3458.5371616616617u,1.5 3459.5137017017014u,1.5 3459.5147017017016u,0 3463.4238618618615u,0 3463.4248618618617u,1.5 3464.401401901902u,1.5 3464.402401901902u,0 3466.356481981982u,0 3466.3574819819823u,1.5 3468.311562062062u,1.5 3468.312562062062u,0 3469.289102102102u,0 3469.290102102102u,1.5 3471.244182182182u,1.5 3471.2451821821824u,0 3472.221722222222u,0 3472.2227222222223u,1.5 3475.1543423423423u,1.5 3475.1553423423425u,0 3476.1318823823826u,0 3476.132882382383u,1.5 3478.0869624624625u,1.5 3478.0879624624627u,0 3480.0420425425427u,0 3480.043042542543u,1.5 3484.9297427427427u,1.5 3484.930742742743u,0 3485.9072827827827u,0 3485.908282782783u,1.5 3486.8848228228226u,1.5 3486.885822822823u,0 3489.8174429429428u,0 3489.818442942943u,1.5 3494.7051431431432u,1.5 3494.7061431431434u,0 3495.682683183183u,0 3495.6836831831833u,1.5 3496.660223223223u,1.5 3496.6612232232233u,0 3498.6153033033033u,0 3498.6163033033035u,1.5 3500.5703833833836u,1.5 3500.571383383384u,0 3501.547923423423u,0 3501.5489234234233u,1.5 3511.3233238238236u,1.5 3511.3243238238238u,0 3512.3008638638635u,0 3512.3018638638637u,1.5 3513.278403903904u,1.5 3513.279403903904u,0 3515.233483983984u,0 3515.2344839839843u,1.5 3521.098724224224u,1.5 3521.0997242242242u,0 3522.076264264264u,0 3522.077264264264u,1.5 3524.0313443443442u,1.5 3524.0323443443444u,0 3525.986424424424u,0 3525.9874244244243u,1.5 3527.9415045045043u,1.5 3527.9425045045045u,0 3528.9190445445447u,0 3528.920044544545u,1.5 3529.8965845845846u,1.5 3529.897584584585u,0 3530.8741246246245u,0 3530.8751246246247u,1.5 3532.8292047047044u,1.5 3532.8302047047046u,0 3538.6944449449447u,0 3538.695444944945u,1.5 3539.671984984985u,1.5 3539.6729849849853u,0 3544.559685185185u,0 3544.5606851851853u,1.5 3545.537225225225u,1.5 3545.5382252252252u,0 3549.4473853853856u,0 3549.448385385386u,1.5 3551.4024654654654u,1.5 3551.4034654654656u,0 3552.3800055055053u,0 3552.3810055055055u,1.5 3553.3575455455457u,1.5 3553.358545545546u,0 3554.3350855855856u,0 3554.336085585586u,1.5 3556.2901656656654u,1.5 3556.2911656656656u,0 3557.2677057057053u,0 3557.2687057057055u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.020646146146u,0 3568.0216461461464u,1.5 3569.975726226226u,1.5 3569.976726226226u,0 3571.9308063063063u,0 3571.9318063063065u,1.5 3572.908346346346u,1.5 3572.9093463463464u,0 3574.863426426426u,0 3574.8644264264262u,1.5 3576.8185065065063u,1.5 3576.8195065065065u,0 3579.7511266266265u,0 3579.7521266266267u,1.5 3586.593906906907u,1.5 3586.594906906907u,0 3587.5714469469467u,0 3587.572446946947u,1.5 3588.548986986987u,1.5 3588.5499869869873u,0 3591.481607107107u,0 3591.482607107107u,1.5 3592.459147147147u,1.5 3592.4601471471474u,0 3593.436687187187u,0 3593.4376871871873u,1.5 3594.414227227227u,1.5 3594.415227227227u,0 3595.391767267267u,0 3595.392767267267u,1.5 3596.3693073073073u,1.5 3596.3703073073075u,0 3597.346847347347u,0 3597.3478473473474u,1.5 3598.3243873873876u,1.5 3598.3253873873878u,0 3599.301927427427u,0 3599.302927427427u,1.5 3602.2345475475477u,1.5 3602.235547547548u,0 3605.1671676676674u,0 3605.1681676676676u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3607.1222477477477u,0 3607.123247747748u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3612.987487987988u,0 3612.9884879879883u,1.5 3613.9650280280275u,1.5 3613.9660280280277u,0 3614.942568068068u,0 3614.943568068068u,1.5 3621.785348348348u,1.5 3621.7863483483484u,0 3623.740428428428u,0 3623.741428428428u,1.5 3624.7179684684684u,1.5 3624.7189684684686u,0 3629.6056686686684u,0 3629.6066686686686u,1.5 3635.4709089089088u,1.5 3635.471908908909u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3637.425988988989u,1.5 3637.4269889889893u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3640.358609109109u,0 3640.359609109109u,1.5 3641.336149149149u,1.5 3641.3371491491494u,0 3644.268769269269u,0 3644.269769269269u,1.5 3645.2463093093093u,1.5 3645.2473093093095u,0 3647.2013893893895u,0 3647.2023893893897u,1.5 3651.1115495495496u,1.5 3651.11254954955u,0 3653.06662962963u,0 3653.06762962963u,1.5 3654.0441696696694u,1.5 3654.0451696696696u,0 3655.0217097097097u,0 3655.02270970971u,1.5 3656.9767897897896u,1.5 3656.9777897897898u,0 3657.95432982983u,0 3657.95532982983u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3669.6848103103102u,0 3669.6858103103104u,1.5 3673.5949704704703u,1.5 3673.5959704704705u,0 3674.5725105105103u,0 3674.5735105105105u,1.5 3675.5500505505506u,1.5 3675.551050550551u,0 3678.4826706706704u,0 3678.4836706706706u,1.5 3679.4602107107107u,1.5 3679.461210710711u,0 3680.4377507507506u,0 3680.438750750751u,1.5 3681.4152907907906u,1.5 3681.4162907907908u,0 3682.392830830831u,0 3682.393830830831u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3689.2356111111108u,1.5 3689.236611111111u,0 3690.213151151151u,0 3690.2141511511513u,1.5 3691.190691191191u,1.5 3691.1916911911912u,0 3693.145771271271u,0 3693.146771271271u,1.5 3697.0559314314314u,1.5 3697.0569314314316u,0 3699.9885515515516u,0 3699.989551551552u,1.5 3700.9660915915915u,1.5 3700.9670915915917u,0 3702.9211716716713u,0 3702.9221716716715u,1.5 3706.831331831832u,1.5 3706.832331831832u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3711.719032032032u,0 3711.720032032032u,1.5 3715.629192192192u,1.5 3715.630192192192u,0 3716.6067322322324u,0 3716.6077322322326u,1.5 3717.584272272272u,1.5 3717.585272272272u,0 3719.539352352352u,0 3719.5403523523523u,1.5 3722.4719724724723u,1.5 3722.4729724724725u,0 3723.4495125125122u,0 3723.4505125125124u,1.5 3724.4270525525526u,1.5 3724.428052552553u,0 3725.4045925925925u,0 3725.4055925925927u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3732.2473728728723u,0 3732.2483728728726u,1.5 3734.2024529529526u,1.5 3734.203452952953u,0 3735.179992992993u,0 3735.180992992993u,1.5 3736.157533033033u,1.5 3736.158533033033u,0 3737.135073073073u,0 3737.136073073073u,1.5 3739.090153153153u,1.5 3739.0911531531533u,0 3740.067693193193u,0 3740.068693193193u,1.5 3741.0452332332334u,1.5 3741.0462332332336u,0 3744.9553933933935u,0 3744.9563933933937u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3753.7532537537536u,1.5 3753.754253753754u,0 3754.730793793794u,0 3754.731793793794u,1.5 3755.708333833834u,1.5 3755.709333833834u,0 3756.685873873874u,0 3756.686873873874u,1.5 3757.6634139139137u,1.5 3757.664413913914u,0 3758.6409539539536u,0 3758.641953953954u,1.5 3759.618493993994u,1.5 3759.619493993994u,0 3760.596034034034u,0 3760.597034034034u,1.5 3761.573574074074u,1.5 3761.574574074074u,0 3764.506194194194u,0 3764.507194194194u,1.5 3772.326514514514u,1.5 3772.3275145145144u,0 3774.2815945945945u,0 3774.2825945945947u,1.5 3775.259134634635u,1.5 3775.260134634635u,0 3776.2366746746743u,0 3776.2376746746745u,1.5 3778.1917547547546u,1.5 3778.192754754755u,0 3779.169294794795u,0 3779.170294794795u,1.5 3780.146834834835u,1.5 3780.147834834835u,0 3781.124374874875u,0 3781.125374874875u,1.5 3783.0794549549546u,1.5 3783.080454954955u,0 3786.012075075075u,0 3786.013075075075u,1.5 3787.967155155155u,1.5 3787.9681551551553u,0 3788.944695195195u,0 3788.945695195195u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3793.8323953953955u,0 3793.8333953953957u,1.5 3794.8099354354354u,1.5 3794.8109354354356u,0 3798.7200955955955u,0 3798.7210955955957u,1.5 3802.6302557557556u,1.5 3802.631255755756u,0 3803.607795795796u,0 3803.608795795796u,1.5 3804.585335835836u,1.5 3804.586335835836u,0 3806.5404159159157u,0 3806.541415915916u,1.5 3808.495495995996u,1.5 3808.496495995996u,0 3809.473036036036u,0 3809.474036036036u,1.5 3812.405656156156u,1.5 3812.4066561561563u,0 3813.383196196196u,0 3813.384196196196u,1.5 3814.3607362362363u,1.5 3814.3617362362365u,0 3815.338276276276u,0 3815.339276276276u,1.5 3821.203516516516u,1.5 3821.2045165165164u,0 3822.1810565565565u,0 3822.1820565565567u,1.5 3825.1136766766763u,1.5 3825.1146766766765u,0 3826.0912167167166u,0 3826.092216716717u,1.5 3828.046296796797u,1.5 3828.047296796797u,0 3831.9564569569566u,0 3831.957456956957u,1.5 3832.933996996997u,1.5 3832.934996996997u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3836.844157157157u,0 3836.8451571571572u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 3844.6644774774772u,0 3844.6654774774775u,1.5 3847.5970975975974u,1.5 3847.5980975975976u,0 3848.574637637638u,0 3848.575637637638u,1.5 3850.5297177177176u,1.5 3850.530717717718u,0 3851.5072577577575u,0 3851.5082577577577u,1.5 3852.484797797798u,1.5 3852.485797797798u,0 3855.4174179179176u,0 3855.418417917918u,1.5 3856.394957957958u,1.5 3856.395957957958u,0 3859.3275780780777u,0 3859.328578078078u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3870.080518518518u,0 3870.0815185185184u,1.5 3873.013138638639u,1.5 3873.014138638639u,0 3873.9906786786783u,0 3873.9916786786785u,1.5 3876.923298798799u,1.5 3876.924298798799u,0 3877.900838838839u,0 3877.901838838839u,1.5 3879.8559189189186u,1.5 3879.856918918919u,0 3888.653779279279u,0 3888.6547792792794u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3895.4965595595595u,1.5 3895.4975595595597u,0 3902.33933983984u,0 3902.34033983984u,1.5 3903.31687987988u,1.5 3903.3178798798804u,0 3904.2944199199196u,0 3904.29541991992u,1.5 3913.09228028028u,1.5 3913.0932802802804u,0 3914.06982032032u,0 3914.0708203203203u,1.5 3915.0473603603605u,1.5 3915.0483603603607u,0 3917.00244044044u,0 3917.00344044044u,1.5 3917.9799804804807u,1.5 3917.980980480481u,0 3919.935060560561u,0 3919.936060560561u,1.5 3920.9126006006004u,1.5 3920.9136006006006u,0 3923.8452207207206u,0 3923.846220720721u,1.5 3925.800300800801u,1.5 3925.801300800801u,0 3926.7778408408403u,0 3926.7788408408405u,1.5 3928.7329209209206u,1.5 3928.733920920921u,0 3929.710460960961u,0 3929.711460960961u,1.5 3933.6206211211206u,1.5 3933.621621121121u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3938.508321321321u,0 3938.5093213213213u,1.5 3939.4858613613615u,1.5 3939.4868613613617u,0 3940.4634014014014u,0 3940.4644014014016u,1.5 3941.440941441441u,1.5 3941.441941441441u,0 3943.396021521521u,0 3943.3970215215213u,1.5 3944.373561561562u,1.5 3944.374561561562u,0 3947.3061816816817u,0 3947.307181681682u,1.5 3948.2837217217216u,1.5 3948.284721721722u,0 3949.261261761762u,0 3949.262261761762u,1.5 3950.238801801802u,1.5 3950.239801801802u,0 3952.193881881882u,0 3952.1948818818823u,1.5 3953.1714219219216u,1.5 3953.172421921922u,0 3954.1489619619624u,0 3954.1499619619626u,1.5 3956.104042042042u,1.5 3956.105042042042u,0 3957.081582082082u,0 3957.0825820820824u,1.5 3960.014202202202u,1.5 3960.015202202202u,0 3961.969282282282u,0 3961.9702822822824u,1.5 3962.946822322322u,1.5 3962.9478223223223u,0 3963.9243623623624u,0 3963.9253623623626u,1.5 3965.879442442442u,1.5 3965.880442442442u,0 3966.8569824824826u,0 3966.857982482483u,1.5 3967.834522522522u,1.5 3967.8355225225223u,0 3969.7896026026024u,0 3969.7906026026026u,1.5 3972.7222227227226u,1.5 3972.7232227227228u,0 3973.699762762763u,0 3973.700762762763u,1.5 3974.677302802803u,1.5 3974.678302802803u,0 3975.6548428428423u,0 3975.6558428428425u,1.5 3977.6099229229226u,1.5 3977.610922922923u,0 3980.5425430430428u,0 3980.543543043043u,1.5 3981.520083083083u,1.5 3981.5210830830833u,0 3982.4976231231226u,0 3982.498623123123u,1.5 3983.4751631631634u,1.5 3983.4761631631636u,0 3989.3404034034033u,0 3989.3414034034035u,1.5 3991.2954834834836u,1.5 3991.296483483484u,0 3998.138263763764u,0 3998.139263763764u,1.5 3999.115803803804u,1.5 3999.116803803804u,0 4000.0933438438433u,0 4000.0943438438435u,1.5 4001.070883883884u,1.5 4001.0718838838843u,0 4013.7789044044043u,0 4013.7799044044045u,1.5 4014.756444444444u,1.5 4014.757444444444u,0 4016.711524524524u,0 4016.7125245245243u,1.5 4018.6666046046043u,1.5 4018.6676046046045u,0 4020.6216846846846u,0 4020.622684684685u,1.5 4021.5992247247245u,1.5 4021.6002247247247u,0 4024.5318448448443u,0 4024.5328448448445u,1.5 4026.4869249249246u,1.5 4026.4879249249248u,0 4027.4644649649654u,0 4027.4654649649656u,1.5 4028.442005005005u,1.5 4028.443005005005u,0 4029.4195450450447u,0 4029.420545045045u,1.5 4030.397085085085u,1.5 4030.3980850850853u,0 4031.374625125125u,0 4031.375625125125u,1.5 4033.329705205205u,1.5 4033.330705205205u,0 4035.284785285285u,0 4035.2857852852853u,1.5 4037.2398653653654u,1.5 4037.2408653653656u,0 4038.2174054054053u,0 4038.2184054054055u,1.5 4039.194945445445u,1.5 4039.195945445445u,0 4040.1724854854856u,0 4040.173485485486u,1.5 4043.1051056056053u,1.5 4043.1061056056055u,0 4045.0601856856856u,0 4045.061185685686u,1.5 4047.015265765766u,1.5 4047.016265765766u,0 4048.9703458458453u,0 4048.9713458458455u,1.5 4049.947885885886u,1.5 4049.9488858858863u,0 4051.9029659659664u,0 4051.9039659659666u,1.5 4052.880506006006u,1.5 4052.881506006006u,0 4057.768206206206u,0 4057.769206206206u,1.5 4058.7457462462457u,1.5 4058.746746246246u,0 4061.6783663663664u,0 4061.6793663663666u,1.5 4062.6559064064063u,1.5 4062.6569064064065u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4065.588526526526u,1.5 4065.5895265265262u,0 4066.566066566567u,0 4066.567066566567u,1.5 4067.5436066066063u,1.5 4067.5446066066065u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4073.4088468468462u,1.5 4073.4098468468464u,0 4074.386386886887u,0 4074.3873868868873u,1.5 4075.3639269269265u,1.5 4075.3649269269267u,0 4076.3414669669673u,0 4076.3424669669675u,1.5 4077.319007007007u,1.5 4077.320007007007u,0 4078.2965470470467u,0 4078.297547047047u,1.5 4079.274087087087u,1.5 4079.2750870870873u,0 4080.251627127127u,0 4080.252627127127u,1.5 4081.2291671671674u,1.5 4081.2301671671676u,0 4084.161787287287u,0 4084.1627872872873u,1.5 4085.139327327327u,1.5 4085.140327327327u,0 4086.1168673673674u,0 4086.1178673673676u,1.5 4087.0944074074073u,1.5 4087.0954074074075u,0 4089.0494874874876u,0 4089.0504874874878u,1.5 4092.959647647647u,1.5 4092.9606476476474u,0 4095.892267767768u,0 4095.893267767768u,1.5 4096.869807807808u,1.5 4096.870807807808u,0 4097.847347847847u,0 4097.848347847847u,1.5 4098.824887887888u,1.5 4098.825887887888u,0 4101.757508008008u,0 4101.758508008008u,1.5 4102.735048048047u,1.5 4102.736048048047u,0 4104.690128128128u,0 4104.691128128128u,1.5 4105.667668168168u,1.5 4105.668668168169u,0 4106.645208208208u,0 4106.646208208208u,1.5 4112.510448448448u,1.5 4112.511448448448u,0 4113.487988488489u,0 4113.488988488489u,1.5 4114.465528528528u,1.5 4114.466528528528u,0 4115.443068568568u,0 4115.444068568569u,1.5 4116.420608608609u,1.5 4116.421608608609u,0 4119.353228728728u,0 4119.354228728728u,1.5 4120.330768768769u,1.5 4120.3317687687695u,0 4122.285848848848u,0 4122.286848848848u,1.5 4124.240928928929u,1.5 4124.241928928929u,0 4125.218468968969u,0 4125.2194689689695u,1.5 4127.173549049048u,1.5 4127.174549049048u,0 4128.1510890890895u,0 4128.15208908909u,1.5 4130.106169169169u,1.5 4130.1071691691695u,0 4131.083709209209u,0 4131.084709209209u,1.5 4132.061249249249u,1.5 4132.062249249249u,0 4134.993869369369u,0 4134.99486936937u,1.5 4137.9264894894895u,1.5 4137.92748948949u,0 4138.904029529529u,0 4138.905029529529u,1.5 4140.85910960961u,1.5 4140.86010960961u,0 4141.836649649649u,0 4141.837649649649u,1.5 4142.81418968969u,1.5 4142.81518968969u,0 4144.76926976977u,0 4144.7702697697705u,1.5 4145.74680980981u,1.5 4145.74780980981u,0 4146.724349849849u,0 4146.725349849849u,1.5 4149.65696996997u,1.5 4149.6579699699705u,0 4150.63451001001u,0 4150.63551001001u,1.5 4154.54467017017u,1.5 4154.5456701701705u,0 4155.52221021021u,0 4155.52321021021u,1.5 4156.49975025025u,1.5 4156.50075025025u,0 4161.38745045045u,0 4161.38845045045u,1.5 4166.27515065065u,1.5 4166.27615065065u,0 4167.2526906906905u,0 4167.253690690691u,1.5 4168.23023073073u,1.5 4168.23123073073u,0 4170.185310810811u,0 4170.186310810811u,1.5 4171.16285085085u,1.5 4171.16385085085u,0 4172.140390890891u,0 4172.141390890891u,1.5 4173.117930930931u,1.5 4173.118930930931u,0 4174.095470970971u,0 4174.0964709709715u,1.5 4178.005631131131u,1.5 4178.006631131131u,0 4178.983171171171u,0 4178.9841711711715u,1.5 4179.960711211211u,1.5 4179.961711211211u,0 4182.893331331331u,0 4182.894331331331u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4190.713651651651u,1.5 4190.714651651651u,0 4192.668731731731u,0 4192.669731731731u,1.5 4194.623811811812u,1.5 4194.624811811812u,0 4197.556431931932u,0 4197.557431931932u,1.5 4198.533971971972u,1.5 4198.5349719719725u,0 4199.511512012012u,0 4199.512512012012u,1.5 4201.4665920920925u,1.5 4201.467592092093u,0 4202.444132132132u,0 4202.445132132132u,1.5 4203.421672172172u,1.5 4203.4226721721725u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4210.264452452452u,0 4210.265452452452u,1.5 4213.197072572572u,1.5 4213.1980725725725u,0 4216.1296926926925u,0 4216.130692692693u,1.5 4217.107232732732u,1.5 4217.108232732732u,0 4219.062312812813u,0 4219.063312812813u,1.5 4222.972472972973u,1.5 4222.9734729729735u,0 4223.950013013013u,0 4223.951013013013u,1.5 4226.882633133133u,1.5 4226.883633133133u,0 4229.815253253253u,0 4229.816253253253u,1.5 4234.702953453453u,1.5 4234.703953453453u,0 4236.658033533533u,0 4236.659033533533u,1.5 4239.590653653653u,1.5 4239.591653653653u,0 4240.5681936936935u,0 4240.569193693694u,1.5 4244.478353853853u,1.5 4244.479353853853u,0 4245.4558938938935u,0 4245.456893893894u,1.5 4246.433433933934u,1.5 4246.434433933934u,0 4251.321134134134u,0 4251.322134134134u,1.5 4254.253754254254u,1.5 4254.254754254254u,0 4255.2312942942945u,0 4255.232294294295u,1.5 4256.208834334334u,1.5 4256.209834334334u,0 4260.1189944944945u,0 4260.119994494495u,1.5 4261.096534534534u,1.5 4261.097534534534u,0 4262.074074574574u,0 4262.0750745745745u,1.5 4265.0066946946945u,1.5 4265.007694694695u,0 4266.961774774775u,0 4266.962774774775u,1.5 4267.939314814815u,1.5 4267.940314814815u,0 4268.916854854855u,0 4268.917854854855u,1.5 4270.871934934935u,1.5 4270.872934934935u,0 4272.827015015015u,0 4272.828015015015u,1.5 4274.782095095095u,1.5 4274.783095095096u,0 4275.759635135135u,0 4275.760635135135u,1.5 4276.737175175175u,1.5 4276.7381751751755u,0 4277.714715215215u,0 4277.715715215215u,1.5 4278.692255255256u,1.5 4278.693255255256u,0 4282.602415415415u,0 4282.603415415415u,1.5 4285.535035535535u,1.5 4285.536035535535u,0 4286.512575575575u,0 4286.5135755755755u,1.5 4288.467655655656u,1.5 4288.468655655656u,0 4289.4451956956955u,0 4289.446195695696u,1.5 4290.422735735735u,1.5 4290.423735735735u,0 4292.377815815816u,0 4292.378815815816u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4294.3328958958955u,0 4294.333895895896u,1.5 4298.243056056056u,1.5 4298.244056056056u,0 4299.220596096096u,0 4299.221596096097u,1.5 4300.198136136136u,1.5 4300.199136136136u,0 4303.130756256257u,0 4303.131756256257u,1.5 4307.040916416417u,1.5 4307.041916416417u,0 4308.018456456457u,0 4308.019456456457u,1.5 4308.995996496496u,1.5 4308.996996496497u,0 4309.973536536536u,0 4309.974536536536u,1.5 4310.951076576576u,1.5 4310.9520765765765u,0 4313.8836966966965u,0 4313.884696696697u,1.5 4317.793856856857u,1.5 4317.794856856857u,0 4318.7713968968965u,0 4318.772396896897u,1.5 4320.726476976977u,1.5 4320.727476976977u,0 4321.704017017017u,0 4321.705017017017u,1.5 4323.659097097097u,1.5 4323.660097097098u,0 4326.591717217217u,0 4326.592717217217u,1.5 4327.569257257258u,1.5 4327.570257257258u,0 4328.546797297297u,0 4328.547797297298u,1.5 4332.456957457458u,1.5 4332.457957457458u,0 4336.367117617618u,0 4336.368117617618u,1.5 4337.344657657658u,1.5 4337.345657657658u,0 4343.2098978978975u,0 4343.210897897898u,1.5 4344.187437937938u,1.5 4344.188437937938u,0 4345.164977977978u,0 4345.165977977978u,1.5 4346.142518018018u,1.5 4346.143518018018u,0 4347.120058058058u,0 4347.121058058058u,1.5 4348.097598098098u,1.5 4348.098598098099u,0 4351.030218218218u,0 4351.031218218218u,1.5 4354.940378378378u,1.5 4354.941378378378u,0 4355.917918418419u,0 4355.918918418419u,1.5 4357.872998498498u,1.5 4357.873998498499u,0 4358.850538538538u,0 4358.851538538538u,1.5 4359.828078578578u,1.5 4359.829078578578u,0 4361.783158658659u,0 4361.784158658659u,1.5 4362.760698698698u,1.5 4362.761698698699u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4368.625938938939u,1.5 4368.626938938939u,0 4370.581019019019u,0 4370.582019019019u,1.5 4371.558559059059u,1.5 4371.559559059059u,0 4372.536099099099u,0 4372.5370990991u,1.5 4374.491179179179u,1.5 4374.492179179179u,0 4375.468719219219u,0 4375.469719219219u,1.5 4377.423799299299u,1.5 4377.4247992993u,0 4379.378879379379u,0 4379.379879379379u,1.5 4382.311499499499u,1.5 4382.3124994995u,0 4383.289039539539u,0 4383.290039539539u,1.5 4385.24411961962u,1.5 4385.24511961962u,0 4386.22165965966u,0 4386.22265965966u,1.5 4387.199199699699u,1.5 4387.2001996997u,0 4390.13181981982u,0 4390.13281981982u,1.5 4391.10935985986u,1.5 4391.11035985986u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.99706006006u,0 4395.99806006006u,1.5 4402.83984034034u,1.5 4402.84084034034u,0 4403.81738038038u,0 4403.81838038038u,1.5 4404.794920420421u,1.5 4404.795920420421u,0 4405.772460460461u,0 4405.773460460461u,1.5 4406.7500005005u,1.5 4406.751000500501u,0 4411.6377007007u,0 4411.638700700701u,1.5 4412.61524074074u,1.5 4412.61624074074u,0 4414.570320820821u,0 4414.571320820821u,1.5 4416.5254009009u,1.5 4416.526400900901u,0 4417.502940940941u,0 4417.503940940941u,1.5 4418.480480980981u,1.5 4418.481480980981u,0 4419.458021021021u,0 4419.459021021021u,1.5 4420.435561061061u,1.5 4420.436561061061u,0 4421.413101101101u,0 4421.414101101102u,1.5 4423.368181181181u,1.5 4423.369181181181u,0 4424.345721221221u,0 4424.346721221221u,1.5 4425.323261261262u,1.5 4425.324261261262u,0 4426.300801301301u,0 4426.301801301302u,1.5 4427.278341341341u,1.5 4427.279341341341u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4438.031281781782u,0 4438.032281781782u,1.5 4440.963901901901u,1.5 4440.964901901902u,0 4441.941441941942u,0 4441.942441941942u,1.5 4442.918981981982u,1.5 4442.919981981982u,0 4443.896522022022u,0 4443.897522022022u,1.5 4448.784222222222u,1.5 4448.785222222222u,0 4450.739302302302u,0 4450.740302302303u,1.5 4451.716842342342u,1.5 4451.717842342342u,0 4452.694382382382u,0 4452.695382382382u,1.5 4453.6719224224225u,1.5 4453.672922422423u,0 4456.604542542542u,0 4456.605542542542u,1.5 4457.582082582582u,1.5 4457.583082582582u,0 4459.537162662663u,0 4459.538162662663u,1.5 4460.514702702702u,1.5 4460.515702702703u,0 4462.469782782783u,0 4462.470782782783u,1.5 4463.447322822823u,1.5 4463.448322822823u,0 4465.402402902902u,0 4465.403402902903u,1.5 4466.379942942943u,1.5 4466.380942942943u,0 4467.357482982983u,0 4467.358482982983u,1.5 4468.335023023023u,1.5 4468.336023023023u,0 4469.312563063063u,0 4469.313563063063u,1.5 4470.290103103103u,1.5 4470.2911031031035u,0 4471.267643143143u,0 4471.268643143143u,1.5 4472.245183183183u,1.5 4472.246183183183u,0 4473.222723223223u,0 4473.223723223223u,1.5 4476.155343343343u,1.5 4476.156343343343u,0 4478.1104234234235u,0 4478.111423423424u,1.5 4479.087963463464u,1.5 4479.088963463464u,0 4480.065503503503u,0 4480.066503503504u,1.5 4488.863363863864u,1.5 4488.864363863864u,0 4495.706144144144u,0 4495.707144144144u,1.5 4496.683684184184u,1.5 4496.684684184184u,0 4497.661224224224u,0 4497.662224224224u,1.5 4502.5489244244245u,1.5 4502.549924424425u,0 4503.526464464465u,0 4503.527464464465u,1.5 4504.504004504504u,1.5 4504.5050045045045u,0 4506.459084584585u,0 4506.460084584585u,1.5 4516.234484984985u,1.5 4516.235484984985u,0 4517.212025025025u,0 4517.213025025025u,1.5 4519.167105105105u,1.5 4519.1681051051055u,0 4520.144645145145u,0 4520.145645145145u,1.5 4521.122185185185u,1.5 4521.123185185185u,0 4523.077265265266u,0 4523.078265265266u,1.5 4524.054805305305u,1.5 4524.0558053053055u,0 4525.032345345345u,0 4525.033345345345u,1.5 4526.009885385385u,1.5 4526.010885385385u,0 4526.9874254254255u,0 4526.988425425426u,1.5 4528.942505505505u,1.5 4528.9435055055055u,0 4530.897585585586u,0 4530.898585585586u,1.5 4532.852665665666u,1.5 4532.853665665666u,0 4534.807745745745u,0 4534.808745745745u,1.5 4535.785285785786u,1.5 4535.786285785786u,0 4546.538226226226u,0 4546.539226226226u,1.5 4547.515766266267u,1.5 4547.516766266267u,0 4549.470846346346u,0 4549.471846346346u,1.5 4551.4259264264265u,1.5 4551.426926426427u,0 4552.403466466467u,0 4552.404466466467u,1.5 4556.3136266266265u,1.5 4556.314626626627u,0 4557.291166666667u,0 4557.292166666667u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4566.0890270270265u,0 4566.090027027027u,1.5 4567.066567067067u,1.5 4567.067567067067u,0 4571.954267267268u,0 4571.955267267268u,1.5 4572.931807307307u,1.5 4572.9328073073075u,0 4575.8644274274275u,0 4575.865427427428u,1.5 4576.841967467468u,1.5 4576.842967467468u,0 4577.819507507507u,0 4577.8205075075075u,1.5 4578.797047547547u,1.5 4578.798047547547u,0 4579.774587587588u,0 4579.775587587588u,1.5 4584.662287787788u,1.5 4584.663287787788u,0 4585.6398278278275u,0 4585.640827827828u,1.5 4586.617367867868u,1.5 4586.618367867868u,0 4597.370308308308u,0 4597.3713083083085u,1.5 4598.347848348348u,1.5 4598.348848348348u,0 4599.325388388388u,0 4599.326388388388u,1.5 4601.280468468469u,1.5 4601.281468468469u,0 4602.258008508508u,0 4602.2590085085085u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4609.100788788789u,0 4609.101788788789u,1.5 4610.0783288288285u,1.5 4610.079328828829u,0 4613.988488988989u,0 4613.989488988989u,1.5 4614.9660290290285u,1.5 4614.967029029029u,0 4615.943569069069u,0 4615.944569069069u,1.5 4616.921109109109u,1.5 4616.922109109109u,0 4617.898649149149u,0 4617.899649149149u,1.5 4620.83126926927u,1.5 4620.83226926927u,0 4623.763889389389u,0 4623.764889389389u,1.5 4624.741429429429u,1.5 4624.74242942943u,0 4627.674049549549u,0 4627.675049549549u,1.5 4630.60666966967u,1.5 4630.60766966967u,0 4631.584209709709u,0 4631.5852097097095u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4636.471909909909u,0 4636.4729099099095u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4641.35961011011u,0 4641.36061011011u,1.5 4642.33715015015u,1.5 4642.33815015015u,0 4643.31469019019u,0 4643.31569019019u,1.5 4644.2922302302295u,1.5 4644.29323023023u,0 4645.269770270271u,0 4645.270770270271u,1.5 4648.20239039039u,1.5 4648.20339039039u,0 4649.17993043043u,0 4649.180930430431u,1.5 4651.13501051051u,1.5 4651.1360105105105u,0 4656.02271071071u,0 4656.0237107107105u,1.5 4657.977790790791u,1.5 4657.978790790791u,0 4658.9553308308305u,0 4658.956330830831u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4667.753191191191u,0 4667.754191191191u,1.5 4675.573511511511u,1.5 4675.574511511511u,0 4680.461211711711u,0 4680.4622117117115u,1.5 4682.416291791792u,1.5 4682.417291791792u,0 4683.393831831831u,0 4683.394831831832u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4689.259072072072u,0 4689.260072072072u,1.5 4690.236612112112u,1.5 4690.237612112112u,0 4691.214152152152u,0 4691.215152152152u,1.5 4693.1692322322315u,1.5 4693.170232232232u,0 4694.146772272273u,0 4694.147772272273u,1.5 4696.101852352352u,1.5 4696.102852352352u,0 4698.056932432432u,0 4698.057932432433u,1.5 4699.034472472473u,1.5 4699.035472472473u,0 4700.012012512512u,0 4700.013012512512u,1.5 4703.922172672673u,1.5 4703.923172672673u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4712.720033033032u,0 4712.721033033033u,1.5 4715.652653153153u,1.5 4715.653653153153u,0 4717.6077332332325u,0 4717.608733233233u,1.5 4718.585273273274u,1.5 4718.586273273274u,0 4719.562813313313u,0 4719.563813313313u,1.5 4720.540353353353u,1.5 4720.541353353353u,0 4723.472973473474u,0 4723.473973473474u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4731.293293793794u,0 4731.294293793794u,1.5 4732.270833833833u,1.5 4732.271833833834u,0 4735.203453953954u,0 4735.204453953954u,1.5 4739.113614114114u,1.5 4739.114614114114u,0 4740.091154154154u,0 4740.092154154154u,1.5 4741.068694194194u,1.5 4741.069694194194u,0 4742.046234234233u,0 4742.047234234234u,1.5 4743.023774274275u,1.5 4743.024774274275u,0 4744.001314314314u,0 4744.002314314314u,1.5 4744.978854354354u,1.5 4744.979854354354u,0 4745.956394394394u,0 4745.957394394394u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4754.7542547547555u,0 4754.755254754756u,1.5 4755.731794794795u,1.5 4755.732794794795u,0 4756.709334834834u,0 4756.710334834835u,1.5 4759.6419549549555u,1.5 4759.642954954956u,0 4760.619494994995u,0 4760.620494994995u,1.5 4761.597035035034u,1.5 4761.598035035035u,0 4763.552115115115u,0 4763.553115115115u,1.5 4764.5296551551555u,1.5 4764.530655155156u,0 4765.507195195195u,0 4765.508195195195u,1.5 4767.462275275276u,1.5 4767.463275275276u,0 4769.4173553553555u,0 4769.418355355356u,1.5 4771.372435435435u,1.5 4771.373435435436u,0 4777.237675675676u,0 4777.238675675676u,1.5 4782.125375875876u,1.5 4782.126375875876u,0 4783.102915915916u,0 4783.103915915916u,1.5 4784.0804559559565u,1.5 4784.081455955957u,0 4787.990616116116u,0 4787.991616116116u,1.5 4793.8558563563565u,1.5 4793.856856356357u,0 4796.788476476477u,0 4796.789476476477u,1.5 4797.766016516516u,1.5 4797.767016516516u,0 4799.721096596597u,0 4799.722096596597u,1.5 4802.653716716716u,1.5 4802.654716716716u,0 4803.6312567567575u,0 4803.632256756758u,1.5 4807.541416916917u,1.5 4807.542416916917u,0 4809.496496996997u,0 4809.497496996997u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4819.271897397397u,0 4819.272897397397u,1.5 4820.249437437437u,1.5 4820.2504374374375u,0 4822.204517517517u,0 4822.205517517517u,1.5 4824.159597597598u,1.5 4824.160597597598u,0 4826.114677677678u,0 4826.115677677678u,1.5 4828.069757757758u,1.5 4828.070757757759u,0 4831.002377877878u,0 4831.003377877878u,1.5 4831.979917917918u,1.5 4831.980917917918u,0 4832.9574579579585u,0 4832.958457957959u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4840.777778278279u,0 4840.778778278279u,1.5 4842.7328583583585u,1.5 4842.733858358359u,0 4844.687938438438u,0 4844.6889384384385u,1.5 4848.598098598599u,1.5 4848.599098598599u,0 4849.575638638638u,0 4849.5766386386385u,1.5 4852.508258758759u,1.5 4852.50925875876u,0 4854.463338838838u,0 4854.464338838839u,1.5 4855.440878878879u,1.5 4855.441878878879u,0 4857.395958958959u,0 4857.39695895896u,1.5 4863.261199199199u,1.5 4863.262199199199u,0 4864.238739239238u,0 4864.239739239239u,1.5 4866.193819319319u,1.5 4866.194819319319u,0 4869.126439439439u,0 4869.1274394394395u,1.5 4870.10397947948u,1.5 4870.10497947948u,0 4871.081519519519u,0 4871.082519519519u,1.5 4872.0590595595595u,1.5 4872.06005955956u,0 4874.014139639639u,0 4874.0151396396395u,1.5 4875.969219719719u,1.5 4875.970219719719u,0 4876.94675975976u,0 4876.947759759761u,1.5 4877.9242997998u,1.5 4877.9252997998u,0 4878.901839839839u,0 4878.9028398398395u,1.5 4879.87937987988u,1.5 4879.88037987988u,0 4880.85691991992u,0 4880.85791991992u,1.5 4881.83445995996u,1.5 4881.835459959961u,0 4883.789540040039u,0 4883.79054004004u,1.5 4884.76708008008u,1.5 4884.76808008008u,0 4886.7221601601605u,0 4886.723160160161u,1.5 4888.677240240239u,1.5 4888.67824024024u,0 4889.654780280281u,0 4889.655780280281u,1.5 4891.6098603603605u,1.5 4891.610860360361u,0 4892.5874004004u,0 4892.5884004004u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4894.542480480481u,0 4894.543480480481u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4898.45264064064u,0 4898.4536406406405u,1.5 4899.430180680681u,1.5 4899.431180680681u,0 4900.40772072072u,0 4900.40872072072u,1.5 4901.385260760761u,1.5 4901.386260760762u,0 4903.34034084084u,0 4903.3413408408405u,1.5 4904.317880880881u,1.5 4904.318880880881u,0 4905.295420920921u,0 4905.296420920921u,1.5 4912.138201201201u,1.5 4912.139201201201u,0 4913.11574124124u,0 4913.116741241241u,1.5 4914.093281281282u,1.5 4914.094281281282u,0 4915.070821321321u,0 4915.071821321321u,1.5 4918.003441441441u,1.5 4918.0044414414415u,0 4919.958521521521u,0 4919.959521521521u,1.5 4920.9360615615615u,1.5 4920.937061561562u,0 4921.913601601602u,0 4921.914601601602u,1.5 4922.891141641641u,1.5 4922.8921416416415u,0 4923.868681681682u,0 4923.869681681682u,1.5 4925.823761761762u,1.5 4925.824761761763u,0 4926.801301801802u,0 4926.802301801802u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4938.531782282283u,1.5 4938.532782282283u,0 4940.486862362362u,0 4940.487862362363u,1.5 4941.464402402402u,1.5 4941.465402402402u,0 4945.3745625625625u,0 4945.375562562563u,1.5 4946.352102602603u,1.5 4946.353102602603u,0 4947.329642642642u,0 4947.3306426426425u,1.5 4948.307182682683u,1.5 4948.308182682683u,0 4949.284722722722u,0 4949.285722722722u,1.5 4950.262262762763u,1.5 4950.263262762764u,0 4953.194882882883u,0 4953.195882882883u,1.5 4954.172422922923u,1.5 4954.173422922923u,0 4955.149962962963u,0 4955.150962962964u,1.5 4956.127503003003u,1.5 4956.128503003003u,0 4957.105043043042u,0 4957.1060430430425u,1.5 4965.902903403403u,1.5 4965.903903403403u,0 4966.880443443443u,0 4966.8814434434435u,1.5 4968.835523523523u,1.5 4968.836523523523u,0 4970.790603603604u,0 4970.791603603604u,1.5 4971.768143643643u,1.5 4971.7691436436435u,0 4972.745683683684u,0 4972.746683683684u,1.5 4973.723223723723u,1.5 4973.724223723723u,0 4974.700763763764u,0 4974.701763763765u,1.5 4975.678303803804u,1.5 4975.679303803804u,0 4976.655843843843u,0 4976.6568438438435u,1.5 4977.633383883884u,1.5 4977.634383883884u,0 4979.588463963964u,0 4979.589463963965u,1.5 4980.566004004004u,1.5 4980.567004004004u,0 4981.543544044043u,0 4981.5445440440435u,1.5 4982.521084084084u,1.5 4982.522084084084u,0 4983.498624124124u,0 4983.499624124124u,1.5 4984.476164164164u,1.5 4984.477164164165u,0 4986.431244244243u,0 4986.4322442442435u,1.5 4987.408784284285u,1.5 4987.409784284285u,0 4988.386324324324u,0 4988.387324324324u,1.5 4991.318944444444u,1.5 4991.319944444444u,0 4992.296484484485u,0 4992.297484484485u,1.5 4993.274024524524u,1.5 4993.275024524524u,0 4994.251564564564u,0 4994.252564564565u,1.5 4995.229104604605u,1.5 4995.230104604605u,0 4996.206644644644u,0 4996.2076446446445u,1.5 4998.161724724724u,1.5 4998.162724724724u,0 5007.937125125125u,0 5007.938125125125u,1.5 5009.892205205205u,1.5 5009.893205205205u,0 5014.779905405405u,0 5014.780905405405u,1.5 5015.757445445445u,1.5 5015.758445445445u,0 5016.734985485486u,0 5016.735985485486u,1.5 5017.712525525525u,1.5 5017.713525525525u,0 5021.622685685686u,0 5021.623685685686u,1.5 5022.600225725725u,1.5 5022.601225725725u,0 5024.555305805806u,0 5024.556305805806u,1.5 5025.532845845845u,1.5 5025.5338458458455u,0 5027.487925925926u,0 5027.488925925926u,1.5 5028.465465965966u,1.5 5028.466465965967u,0 5029.443006006006u,0 5029.444006006006u,1.5 5030.420546046045u,1.5 5030.4215460460455u,0 5031.398086086087u,0 5031.399086086087u,1.5 5033.353166166166u,1.5 5033.354166166167u,0 5035.308246246245u,0 5035.3092462462455u,1.5 5039.218406406406u,1.5 5039.219406406406u,0 5040.195946446446u,0 5040.196946446446u,1.5 5043.128566566566u,1.5 5043.129566566567u,0 5044.106106606607u,0 5044.107106606607u,1.5 5046.061186686687u,1.5 5046.062186686687u,0 5047.038726726726u,0 5047.039726726726u,1.5 5049.971346846846u,1.5 5049.972346846846u,0 5050.948886886887u,0 5050.949886886887u,1.5 5052.903966966967u,1.5 5052.904966966968u,0 5057.791667167167u,0 5057.792667167168u,1.5 5058.769207207207u,1.5 5058.770207207207u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5064.634447447447u,0 5064.635447447447u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5068.544607607608u,1.5 5068.545607607608u,0 5069.522147647647u,0 5069.523147647647u,1.5 5076.364927927928u,1.5 5076.365927927928u,0 5078.320008008008u,0 5078.321008008008u,1.5 5079.297548048047u,1.5 5079.298548048047u,0 5083.207708208208u,0 5083.208708208208u,1.5 5084.185248248248u,1.5 5084.186248248248u,0 5086.140328328328u,0 5086.141328328328u,1.5 5087.117868368368u,1.5 5087.118868368369u,0 5088.095408408408u,0 5088.096408408408u,1.5 5090.050488488489u,1.5 5090.051488488489u,0 5093.960648648648u,0 5093.961648648648u,1.5 5096.893268768769u,1.5 5096.8942687687695u,0 5097.870808808809u,0 5097.871808808809u,1.5 5098.848348848848u,1.5 5098.849348848848u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5112.533909409409u,1.5 5112.534909409409u,0 5113.511449449449u,0 5113.512449449449u,1.5 5114.4889894894895u,1.5 5114.48998948949u,0 5115.466529529529u,0 5115.467529529529u,1.5 5116.444069569569u,1.5 5116.44506956957u,0 5120.354229729729u,0 5120.355229729729u,1.5 5121.33176976977u,1.5 5121.3327697697705u,0 5123.286849849849u,0 5123.287849849849u,1.5 5124.26438988989u,1.5 5124.26538988989u,0 5125.24192992993u,0 5125.24292992993u,1.5 5128.174550050049u,1.5 5128.175550050049u,0 5129.1520900900905u,0 5129.153090090091u,1.5 5130.12963013013u,1.5 5130.13063013013u,0 5131.10717017017u,0 5131.1081701701705u,1.5 5132.08471021021u,1.5 5132.08571021021u,0 5135.01733033033u,0 5135.01833033033u,1.5 5135.99487037037u,1.5 5135.9958703703705u,0 5136.97241041041u,0 5136.97341041041u,1.5 5142.83765065065u,1.5 5142.83865065065u,0 5143.8151906906905u,0 5143.816190690691u,1.5 5144.79273073073u,1.5 5144.79373073073u,0 5149.680430930931u,0 5149.681430930931u,1.5 5150.657970970971u,1.5 5150.6589709709715u,0 5152.61305105105u,0 5152.61405105105u,1.5 5153.5905910910915u,1.5 5153.591591091092u,0 5156.523211211211u,0 5156.524211211211u,1.5 5157.500751251251u,1.5 5157.501751251251u,0 5158.4782912912915u,0 5158.479291291292u,1.5 5159.455831331331u,1.5 5159.456831331331u,0 5160.433371371371u,0 5160.4343713713715u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5162.388451451451u,0 5162.389451451451u,1.5 5168.2536916916915u,1.5 5168.254691691692u,0 5170.208771771772u,0 5170.2097717717725u,1.5 5172.163851851851u,1.5 5172.164851851851u,0 5174.118931931932u,0 5174.119931931932u,1.5 5176.074012012012u,1.5 5176.075012012012u,0 5177.051552052051u,0 5177.052552052051u,1.5 5181.939252252252u,1.5 5181.940252252252u,0 5186.826952452452u,0 5186.827952452452u,1.5 5190.737112612613u,1.5 5190.738112612613u,0 5193.669732732732u,0 5193.670732732732u,1.5 5195.624812812813u,1.5 5195.625812812813u,0 5198.557432932933u,0 5198.558432932933u,1.5 5199.534972972973u,1.5 5199.5359729729735u,0 5200.512513013013u,0 5200.513513013013u,1.5 5201.490053053052u,1.5 5201.491053053052u,0 5202.4675930930935u,0 5202.468593093094u,1.5 5203.445133133133u,1.5 5203.446133133133u,0 5208.332833333333u,0 5208.333833333333u,1.5 5213.220533533533u,1.5 5213.221533533533u,0 5218.108233733733u,0 5218.109233733733u,1.5 5220.063313813814u,1.5 5220.064313813814u,0 5221.040853853853u,0 5221.041853853853u,1.5 5222.995933933934u,1.5 5222.996933933934u,0 5223.973473973974u,0 5223.974473973974u,1.5 5225.928554054053u,1.5 5225.929554054053u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5232.771334334334u,0 5232.772334334334u,1.5 5235.703954454454u,1.5 5235.704954454454u,0 5237.659034534534u,0 5237.660034534534u,1.5 5238.636574574574u,1.5 5238.6375745745745u,0 5240.591654654654u,0 5240.592654654654u,1.5 5244.501814814815u,1.5 5244.502814814815u,0 5250.367055055054u,0 5250.368055055054u,1.5 5254.277215215215u,1.5 5254.278215215215u,0 5255.254755255255u,0 5255.255755255255u,1.5 5256.232295295295u,1.5 5256.233295295296u,0 5258.187375375375u,0 5258.1883753753755u,1.5 5261.1199954954955u,1.5 5261.120995495496u,0 5262.097535535535u,0 5262.098535535535u,1.5 5266.0076956956955u,1.5 5266.008695695696u,0 5271.872935935936u,0 5271.873935935936u,1.5 5275.783096096096u,1.5 5275.784096096097u,0 5276.760636136136u,0 5276.761636136136u,1.5 5277.738176176176u,1.5 5277.739176176176u,0 5280.670796296296u,0 5280.671796296297u,1.5 5281.648336336336u,1.5 5281.649336336336u,0 5282.625876376376u,0 5282.6268763763765u,1.5 5283.603416416417u,1.5 5283.604416416417u,0 5285.558496496496u,0 5285.559496496497u,1.5 5287.513576576576u,1.5 5287.5145765765765u,0 5288.491116616617u,0 5288.492116616617u,1.5 5290.4461966966965u,1.5 5290.447196696697u,0 5292.401276776777u,0 5292.402276776777u,1.5 5294.356356856857u,1.5 5294.357356856857u,0 5295.3338968968965u,0 5295.334896896897u,1.5 5296.311436936937u,1.5 5296.312436936937u,0 5297.288976976977u,0 5297.289976976977u,1.5 5300.221597097097u,1.5 5300.222597097098u,0 5302.176677177177u,0 5302.177677177177u,1.5 5303.154217217217u,1.5 5303.155217217217u,0 5304.131757257258u,0 5304.132757257258u,1.5 5305.109297297297u,1.5 5305.110297297298u,0 5306.086837337337u,0 5306.087837337337u,1.5 5307.064377377377u,1.5 5307.065377377377u,0 5308.041917417418u,0 5308.042917417418u,1.5 5309.019457457458u,1.5 5309.020457457458u,0 5312.929617617618u,0 5312.930617617618u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5320.749937937938u,1.5 5320.750937937938u,0 5322.705018018018u,0 5322.706018018018u,1.5 5323.682558058058u,1.5 5323.683558058058u,0 5326.615178178178u,0 5326.616178178178u,1.5 5327.592718218218u,1.5 5327.593718218218u,0 5329.547798298298u,0 5329.548798298299u,1.5 5330.525338338338u,1.5 5330.526338338338u,0 5331.502878378378u,0 5331.503878378378u,1.5 5332.480418418419u,1.5 5332.481418418419u,0 5334.435498498498u,0 5334.436498498499u,1.5 5335.413038538538u,1.5 5335.414038538538u,0 5337.368118618619u,0 5337.369118618619u,1.5 5338.345658658659u,1.5 5338.346658658659u,0 5339.323198698698u,0 5339.324198698699u,1.5 5344.210898898898u,1.5 5344.211898898899u,0 5353.00875925926u,0 5353.00975925926u,1.5 5354.963839339339u,1.5 5354.964839339339u,0 5356.91891941942u,0 5356.91991941942u,1.5 5357.89645945946u,1.5 5357.89745945946u,0 5361.80661961962u,0 5361.80761961962u,1.5 5363.761699699699u,1.5 5363.7626996997u,0 5364.739239739739u,0 5364.740239739739u,1.5 5366.69431981982u,1.5 5366.69531981982u,0 5368.649399899899u,0 5368.6503998999u,1.5 5371.58202002002u,1.5 5371.58302002002u,0 5374.51464014014u,0 5374.51564014014u,1.5 5375.49218018018u,1.5 5375.49318018018u,0 5376.46972022022u,0 5376.47072022022u,1.5 5377.447260260261u,1.5 5377.448260260261u,0 5378.4248003003u,0 5378.425800300301u,1.5 5386.245120620621u,1.5 5386.246120620621u,0 5394.065440940941u,0 5394.066440940941u,1.5 5395.042980980981u,1.5 5395.043980980981u,0 5396.020521021021u,0 5396.021521021021u,1.5 5396.998061061061u,1.5 5396.999061061061u,0 5397.975601101101u,0 5397.976601101102u,1.5 5398.953141141141u,1.5 5398.954141141141u,0 5399.930681181181u,0 5399.931681181181u,1.5 5400.908221221221u,1.5 5400.909221221221u,0 5401.885761261262u,0 5401.886761261262u,1.5 5402.863301301301u,1.5 5402.864301301302u,0 5406.773461461462u,0 5406.774461461462u,1.5 5408.728541541541u,1.5 5408.729541541541u,0 5409.706081581581u,0 5409.707081581581u,1.5 5411.661161661662u,1.5 5411.662161661662u,0 5413.616241741741u,0 5413.617241741741u,1.5 5421.436562062062u,1.5 5421.437562062062u,0 5422.414102102102u,0 5422.4151021021025u,1.5 5424.369182182182u,1.5 5424.370182182182u,0 5425.346722222222u,0 5425.347722222222u,1.5 5426.324262262263u,1.5 5426.325262262263u,0 5429.256882382382u,0 5429.257882382382u,1.5 5431.211962462463u,1.5 5431.212962462463u,0 5432.189502502502u,0 5432.190502502503u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5438.054742742742u,1.5 5438.055742742742u,0 5439.032282782783u,0 5439.033282782783u,1.5 5440.009822822823u,1.5 5440.010822822823u,0 5440.987362862863u,0 5440.988362862863u,1.5 5443.919982982983u,1.5 5443.920982982983u,0 5445.875063063063u,0 5445.876063063063u,1.5 5446.852603103103u,1.5 5446.8536031031035u,0 5447.830143143143u,0 5447.831143143143u,1.5 5448.807683183183u,1.5 5448.808683183183u,0 5450.762763263264u,0 5450.763763263264u,1.5 5451.740303303303u,1.5 5451.7413033033035u,0 5457.605543543543u,0 5457.606543543543u,1.5 5458.583083583583u,1.5 5458.584083583583u,0 5461.515703703703u,0 5461.516703703704u,1.5 5462.493243743743u,1.5 5462.494243743743u,0 5464.448323823824u,0 5464.449323823824u,1.5 5465.425863863864u,1.5 5465.426863863864u,0 5470.313564064064u,0 5470.314564064064u,1.5 5471.291104104104u,1.5 5471.2921041041045u,0 5473.246184184184u,0 5473.247184184184u,1.5 5474.223724224224u,1.5 5474.224724224224u,0 5475.201264264265u,0 5475.202264264265u,1.5 5478.133884384384u,1.5 5478.134884384384u,0 5479.1114244244245u,0 5479.112424424425u,1.5 5480.088964464465u,1.5 5480.089964464465u,0 5482.044044544544u,0 5482.045044544544u,1.5 5483.021584584585u,1.5 5483.022584584585u,0 5485.954204704704u,0 5485.955204704705u,1.5 5486.931744744744u,1.5 5486.932744744744u,0 5487.909284784785u,0 5487.910284784785u,1.5 5488.8868248248245u,1.5 5488.887824824825u,0 5489.864364864865u,0 5489.865364864865u,1.5 5490.841904904904u,1.5 5490.842904904905u,0 5491.819444944945u,0 5491.820444944945u,1.5 5492.796984984985u,1.5 5492.797984984985u,0 5494.752065065065u,0 5494.753065065065u,1.5 5495.729605105105u,1.5 5495.7306051051055u,0 5496.707145145145u,0 5496.708145145145u,1.5 5499.639765265266u,1.5 5499.640765265266u,0 5500.617305305305u,0 5500.6183053053055u,1.5 5503.5499254254255u,1.5 5503.550925425426u,0 5504.527465465466u,0 5504.528465465466u,1.5 5509.415165665666u,1.5 5509.416165665666u,0 5512.347785785786u,0 5512.348785785786u,1.5 5515.280405905905u,1.5 5515.281405905906u,0 5516.257945945946u,0 5516.258945945946u,1.5 5517.235485985986u,1.5 5517.236485985986u,0 5518.213026026026u,0 5518.214026026026u,1.5 5520.168106106106u,1.5 5520.1691061061065u,0 5521.145646146146u,0 5521.146646146146u,1.5 5524.078266266267u,1.5 5524.079266266267u,0 5525.055806306306u,0 5525.0568063063065u,1.5 5526.033346346346u,1.5 5526.034346346346u,0 5527.010886386386u,0 5527.011886386386u,1.5 5527.9884264264265u,1.5 5527.989426426427u,0 5529.943506506506u,0 5529.9445065065065u,1.5 5530.921046546546u,1.5 5530.922046546546u,0 5531.898586586587u,0 5531.899586586587u,1.5 5533.853666666667u,1.5 5533.854666666667u,0 5538.741366866867u,0 5538.742366866867u,1.5 5539.718906906906u,1.5 5539.7199069069065u,0 5540.696446946947u,0 5540.697446946947u,1.5 5541.673986986987u,1.5 5541.674986986987u,0 5542.6515270270265u,0 5542.652527027027u,1.5 5543.629067067067u,1.5 5543.630067067067u,0 5547.539227227227u,0 5547.540227227227u,1.5 5548.516767267268u,1.5 5548.517767267268u,0 5549.494307307307u,0 5549.4953073073075u,1.5 5550.471847347347u,1.5 5550.472847347347u,0 5552.4269274274275u,0 5552.427927427428u,1.5 5557.3146276276275u,1.5 5557.315627627628u,0 5560.247247747748u,0 5560.248247747748u,1.5 5562.2023278278275u,1.5 5562.203327827828u,0 5563.179867867868u,0 5563.180867867868u,1.5 5566.112487987988u,1.5 5566.113487987988u,0 5567.0900280280275u,0 5567.091028028028u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5570.022648148148u,0 5570.023648148148u,1.5 5571.000188188188u,1.5 5571.001188188188u,0 5572.955268268269u,0 5572.956268268269u,1.5 5573.932808308308u,1.5 5573.9338083083085u,0 5575.887888388388u,0 5575.888888388388u,1.5 5577.842968468469u,1.5 5577.843968468469u,0 5578.820508508508u,0 5578.8215085085085u,1.5 5579.798048548548u,1.5 5579.799048548548u,0 5580.775588588589u,0 5580.776588588589u,1.5 5584.685748748749u,1.5 5584.686748748749u,0 5585.663288788789u,0 5585.664288788789u,1.5 5586.6408288288285u,1.5 5586.641828828829u,0 5587.618368868869u,0 5587.619368868869u,1.5 5589.573448948949u,1.5 5589.574448948949u,0 5595.438689189189u,0 5595.439689189189u,1.5 5596.4162292292285u,1.5 5596.417229229229u,0 5597.39376926927u,0 5597.39476926927u,1.5 5600.326389389389u,1.5 5600.327389389389u,0 5601.303929429429u,0 5601.30492942943u,1.5 5605.21408958959u,1.5 5605.21508958959u,0 5608.146709709709u,0 5608.1477097097095u,1.5 5609.12424974975u,1.5 5609.12524974975u,0 5610.10178978979u,0 5610.10278978979u,1.5 5611.0793298298295u,1.5 5611.08032982983u,0 5613.034409909909u,0 5613.0354099099095u,1.5 5614.01194994995u,1.5 5614.01294994995u,0 5614.98948998999u,0 5614.99048998999u,1.5 5615.9670300300295u,1.5 5615.96803003003u,0 5616.94457007007u,0 5616.94557007007u,1.5 5620.8547302302295u,1.5 5620.85573023023u,0 5621.832270270271u,0 5621.833270270271u,1.5 5623.78735035035u,1.5 5623.78835035035u,0 5628.67505055055u,0 5628.67605055055u,1.5 5629.652590590591u,1.5 5629.653590590591u,0 5630.63013063063u,0 5630.631130630631u,1.5 5632.58521071071u,1.5 5632.5862107107105u,0 5634.540290790791u,0 5634.541290790791u,1.5 5636.495370870871u,1.5 5636.496370870871u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5638.450450950951u,1.5 5638.451450950951u,0 5641.383071071071u,0 5641.384071071071u,1.5 5642.360611111111u,1.5 5642.361611111111u,0 5644.315691191191u,0 5644.316691191191u,1.5 5648.225851351351u,1.5 5648.226851351351u,0 5649.203391391391u,0 5649.204391391391u,1.5 5650.180931431431u,1.5 5650.181931431432u,0 5651.158471471472u,0 5651.159471471472u,1.5 5652.136011511511u,1.5 5652.137011511511u,0 5653.113551551551u,0 5653.114551551551u,1.5 5655.068631631631u,1.5 5655.069631631632u,0 5657.023711711711u,0 5657.0247117117115u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5664.8440320320315u,0 5664.845032032032u,1.5 5665.821572072072u,1.5 5665.822572072072u,0 5666.799112112112u,0 5666.800112112112u,1.5 5667.776652152152u,1.5 5667.777652152152u,0 5669.7317322322315u,0 5669.732732232232u,1.5 5675.596972472473u,1.5 5675.597972472473u,0 5676.574512512512u,0 5676.575512512512u,1.5 5678.529592592593u,1.5 5678.530592592593u,0 5679.507132632632u,0 5679.508132632633u,1.5 5680.484672672673u,1.5 5680.485672672673u,0 5683.417292792793u,0 5683.418292792793u,1.5 5684.394832832832u,1.5 5684.395832832833u,0 5688.304992992993u,0 5688.305992992993u,1.5 5689.282533033032u,1.5 5689.283533033033u,0 5690.260073073073u,0 5690.261073073073u,1.5 5691.237613113113u,1.5 5691.238613113113u,0 5692.215153153153u,0 5692.216153153153u,1.5 5695.147773273274u,1.5 5695.148773273274u,0 5696.125313313313u,0 5696.126313313313u,1.5 5699.057933433433u,1.5 5699.058933433434u,0 5700.035473473474u,0 5700.036473473474u,1.5 5701.013013513513u,1.5 5701.014013513513u,0 5702.968093593594u,0 5702.969093593594u,1.5 5703.945633633633u,1.5 5703.946633633634u,0 5704.923173673674u,0 5704.924173673674u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5711.765953953954u,0 5711.766953953954u,1.5 5713.721034034033u,1.5 5713.722034034034u,0 5716.653654154154u,0 5716.654654154154u,1.5 5718.608734234233u,1.5 5718.609734234234u,0 5722.518894394394u,0 5722.519894394394u,1.5 5723.496434434434u,1.5 5723.497434434435u,0 5725.451514514514u,0 5725.452514514514u,1.5 5726.429054554554u,1.5 5726.430054554554u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5734.249374874875u,0 5734.250374874875u,1.5 5740.114615115115u,1.5 5740.115615115115u,0 5744.024775275276u,0 5744.025775275276u,1.5 5745.002315315315u,1.5 5745.003315315315u,0 5746.957395395395u,0 5746.958395395395u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 5755.7552557557565u,0 5755.756255755757u,1.5 5757.710335835835u,1.5 5757.711335835836u,0 5759.665415915916u,0 5759.666415915916u,1.5 5760.6429559559565u,1.5 5760.643955955957u,0 5761.620495995996u,0 5761.621495995996u,1.5 5762.598036036035u,1.5 5762.599036036036u,0 5764.553116116116u,0 5764.554116116116u,1.5 5766.508196196196u,1.5 5766.509196196196u,0 5767.485736236235u,0 5767.486736236236u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5772.373436436436u,1.5 5772.374436436437u,0 5775.3060565565565u,0 5775.307056556557u,1.5 5776.283596596597u,1.5 5776.284596596597u,0 5777.261136636636u,0 5777.262136636637u,1.5 5778.238676676677u,1.5 5778.239676676677u,0 5779.216216716716u,0 5779.217216716716u,1.5 5780.1937567567575u,1.5 5780.194756756758u,0 5782.148836836836u,0 5782.149836836837u,1.5 5783.126376876877u,1.5 5783.127376876877u,0 5785.0814569569575u,0 5785.082456956958u,1.5 5786.058996996997u,1.5 5786.059996996997u,0 5787.036537037036u,0 5787.037537037037u,1.5 5788.014077077077u,1.5 5788.015077077077u,0 5792.901777277278u,0 5792.902777277278u,1.5 5793.879317317317u,1.5 5793.880317317317u,0 5794.8568573573575u,0 5794.857857357358u,1.5 5795.834397397397u,1.5 5795.835397397397u,0 5798.767017517517u,0 5798.768017517517u,1.5 5799.7445575575575u,1.5 5799.745557557558u,0 5801.699637637637u,0 5801.700637637638u,1.5 5802.677177677678u,1.5 5802.678177677678u,0 5809.5199579579585u,0 5809.520957957959u,1.5 5813.430118118118u,1.5 5813.431118118118u,0 5815.385198198198u,0 5815.386198198198u,1.5 5817.340278278279u,1.5 5817.341278278279u,0 5821.250438438438u,0 5821.2514384384385u,1.5 5822.227978478479u,1.5 5822.228978478479u,0 5823.205518518518u,0 5823.206518518518u,1.5 5825.160598598599u,1.5 5825.161598598599u,0 5827.115678678679u,0 5827.116678678679u,1.5 5829.070758758759u,1.5 5829.07175875876u,0 5830.048298798799u,0 5830.049298798799u,1.5 5831.025838838838u,1.5 5831.026838838839u,0 5833.958458958959u,0 5833.95945895896u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5838.8461591591595u,0 5838.84715915916u,1.5 5840.801239239238u,1.5 5840.802239239239u,0 5842.756319319319u,0 5842.757319319319u,1.5 5843.7338593593595u,1.5 5843.73485935936u,0 5845.688939439439u,0 5845.6899394394395u,1.5 5849.5990995996u,1.5 5849.6000995996u,0 5851.55417967968u,0 5851.55517967968u,1.5 5852.531719719719u,1.5 5852.532719719719u,0 5856.44187987988u,0 5856.44287987988u,1.5 5858.39695995996u,1.5 5858.397959959961u,0 5860.352040040039u,0 5860.35304004004u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5871.104980480481u,0 5871.105980480481u,1.5 5872.08252052052u,1.5 5872.08352052052u,0 5873.0600605605605u,0 5873.061060560561u,1.5 5876.97022072072u,1.5 5876.97122072072u,0 5877.947760760761u,0 5877.948760760762u,1.5 5878.925300800801u,1.5 5878.926300800801u,0 5880.880380880881u,0 5880.881380880881u,1.5 5882.835460960961u,1.5 5882.836460960962u,0 5883.813001001001u,0 5883.814001001001u,1.5 5884.79054104104u,1.5 5884.791541041041u,0 5885.768081081081u,0 5885.769081081081u,1.5 5886.745621121121u,1.5 5886.746621121121u,0 5889.67824124124u,0 5889.679241241241u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5899.453641641641u,0 5899.4546416416415u,1.5 5901.408721721721u,1.5 5901.409721721721u,0 5903.363801801802u,0 5903.364801801802u,1.5 5906.296421921922u,1.5 5906.297421921922u,0 5907.273961961962u,0 5907.274961961963u,1.5 5908.251502002002u,1.5 5908.252502002002u,0 5911.184122122122u,0 5911.185122122122u,1.5 5912.161662162162u,1.5 5912.162662162163u,0 5920.959522522522u,0 5920.960522522522u,1.5 5921.9370625625625u,1.5 5921.938062562563u,0 5922.914602602603u,0 5922.915602602603u,1.5 5923.892142642642u,1.5 5923.8931426426425u,0 5924.869682682683u,0 5924.870682682683u,1.5 5925.847222722722u,1.5 5925.848222722722u,0 5926.824762762763u,0 5926.825762762764u,1.5 5931.712462962963u,1.5 5931.713462962964u,0 5933.667543043042u,0 5933.6685430430425u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5936.600163163163u,0 5936.601163163164u,1.5 5938.555243243242u,1.5 5938.5562432432425u,0 5946.375563563563u,0 5946.376563563564u,1.5 5947.353103603604u,1.5 5947.354103603604u,0 5948.330643643643u,0 5948.3316436436435u,1.5 5949.308183683684u,1.5 5949.309183683684u,0 5950.285723723723u,0 5950.286723723723u,1.5 5951.263263763764u,1.5 5951.264263763765u,0 5952.240803803804u,0 5952.241803803804u,1.5 5953.218343843843u,1.5 5953.2193438438435u,0 5954.195883883884u,0 5954.196883883884u,1.5 5957.128504004004u,1.5 5957.129504004004u,0 5959.083584084084u,0 5959.084584084084u,1.5 5960.061124124124u,1.5 5960.062124124124u,0 5961.038664164164u,0 5961.039664164165u,1.5 5962.993744244243u,1.5 5962.9947442442435u,0 5964.948824324324u,0 5964.949824324324u,1.5 5968.858984484485u,1.5 5968.859984484485u,0 5970.814064564564u,0 5970.815064564565u,1.5 5971.791604604605u,1.5 5971.792604604605u,0 5972.769144644644u,0 5972.7701446446445u,1.5 5973.746684684685u,1.5 5973.747684684685u,0 5979.611924924925u,0 5979.612924924925u,1.5 5980.589464964965u,1.5 5980.590464964966u,0 5983.522085085086u,0 5983.523085085086u,1.5 5984.499625125125u,1.5 5984.500625125125u,0 5986.454705205205u,0 5986.455705205205u,1.5 5987.432245245244u,1.5 5987.4332452452445u,0 6006.005506006006u,0 6006.006506006006u,1.5 6006.983046046045u,1.5 6006.9840460460455u,0 6012.848286286287u,0 6012.849286286287u,1.5 6013.825826326326u,1.5 6013.826826326326u,0 6017.735986486487u,0 6017.736986486487u,1.5 6018.713526526526u,1.5 6018.714526526526u,0 6023.601226726726u,0 6023.602226726726u,1.5 6024.578766766767u,1.5 6024.5797667667675u,0 6028.488926926927u,0 6028.489926926927u,1.5 6029.466466966967u,1.5 6029.467466966968u,0 6030.444007007007u,0 6030.445007007007u,1.5 6032.3990870870875u,1.5 6032.400087087088u,0 6033.376627127127u,0 6033.377627127127u,1.5 6036.309247247247u,1.5 6036.310247247247u,0 6038.264327327327u,0 6038.265327327327u,1.5 6044.129567567567u,1.5 6044.130567567568u,0 6045.107107607608u,0 6045.108107607608u,1.5 6049.994807807808u,1.5 6049.995807807808u,0 6054.882508008008u,0 6054.883508008008u,1.5 6057.815128128128u,1.5 6057.816128128128u,0 6059.770208208208u,0 6059.771208208208u,1.5 6060.747748248248u,1.5 6060.748748248248u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6068.568068568568u,1.5 6068.569068568569u,0 6073.455768768769u,0 6073.4567687687695u,1.5 6074.433308808809u,1.5 6074.434308808809u,0 6075.410848848848u,0 6075.411848848848u,1.5 6076.388388888889u,1.5 6076.389388888889u,0 6077.365928928929u,0 6077.366928928929u,1.5 6078.343468968969u,1.5 6078.3444689689695u,0 6079.321009009009u,0 6079.322009009009u,1.5 6080.298549049048u,1.5 6080.299549049048u,0 6087.141329329329u,0 6087.142329329329u,1.5 6088.118869369369u,1.5 6088.11986936937u,0 6090.073949449449u,0 6090.074949449449u,1.5 6095.93918968969u,1.5 6095.94018968969u,0 6096.916729729729u,0 6096.917729729729u,1.5 6097.89426976977u,1.5 6097.8952697697705u,0 6100.82688988989u,0 6100.82788988989u,1.5 6102.78196996997u,1.5 6102.7829699699705u,0 6103.75951001001u,0 6103.76051001001u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6106.69213013013u,0 6106.69313013013u,1.5 6107.66967017017u,1.5 6107.6706701701705u,0 6108.64721021021u,0 6108.64821021021u,1.5 6113.53491041041u,1.5 6113.53591041041u,0 6117.44507057057u,0 6117.446070570571u,1.5 6130.1530910910915u,1.5 6130.154091091092u,0 6136.018331331331u,0 6136.019331331331u,1.5 6137.973411411411u,1.5 6137.974411411411u,0 6141.883571571571u,0 6141.8845715715715u,1.5 6143.838651651651u,1.5 6143.839651651651u,0 6147.748811811812u,0 6147.749811811812u,1.5 6148.726351851851u,1.5 6148.727351851851u,0 6153.614052052051u,0 6153.615052052051u,1.5 6155.569132132132u,1.5 6155.570132132132u,0 6156.546672172172u,0 6156.5476721721725u,1.5 6157.524212212212u,1.5 6157.525212212212u,0 6158.501752252252u,0 6158.502752252252u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6162.411912412412u,0 6162.412912412412u,1.5 6168.277152652652u,1.5 6168.278152652652u,0 6171.209772772773u,0 6171.210772772773u,1.5 6173.164852852852u,1.5 6173.165852852852u,0 6175.119932932933u,0 6175.120932932933u,1.5 6176.097472972973u,1.5 6176.0984729729735u,0 6177.075013013013u,0 6177.076013013013u,1.5 6178.052553053052u,1.5 6178.053553053052u,0 6179.0300930930935u,0 6179.031093093094u,1.5 6180.985173173173u,1.5 6180.9861731731735u,0 6181.962713213213u,0 6181.963713213213u,1.5 6182.940253253253u,1.5 6182.941253253253u,0 6184.895333333333u,0 6184.896333333333u,1.5 6185.872873373373u,1.5 6185.8738733733735u,0 6186.850413413413u,0 6186.851413413413u,1.5 6190.760573573573u,1.5 6190.7615735735735u,0 6191.738113613614u,0 6191.739113613614u,1.5 6192.715653653653u,1.5 6192.716653653653u,0 6197.603353853853u,0 6197.604353853853u,1.5 6200.535973973974u,1.5 6200.536973973974u,0 6202.491054054053u,0 6202.492054054053u,1.5 6203.468594094094u,1.5 6203.469594094095u,0 6208.3562942942945u,0 6208.357294294295u,1.5 6213.2439944944945u,1.5 6213.244994494495u,0 6215.199074574574u,0 6215.2000745745745u,1.5 6216.176614614615u,1.5 6216.177614614615u,0 6219.109234734734u,0 6219.110234734734u,1.5 6220.086774774775u,1.5 6220.087774774775u,0 6222.041854854854u,0 6222.042854854854u,1.5 6223.0193948948945u,1.5 6223.020394894895u,0 6223.996934934935u,0 6223.997934934935u,1.5 6224.974474974975u,1.5 6224.975474974975u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6233.772335335335u,0 6233.773335335335u,1.5 6235.727415415415u,1.5 6235.728415415415u,0 6238.660035535535u,0 6238.661035535535u,1.5 6244.525275775776u,1.5 6244.526275775776u,0 6245.502815815816u,0 6245.503815815816u,1.5 6246.480355855855u,1.5 6246.481355855855u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6254.300676176176u,0 6254.301676176176u,1.5 6258.210836336336u,1.5 6258.211836336336u,0 6260.165916416417u,0 6260.166916416417u,1.5 6261.143456456457u,1.5 6261.144456456457u,0 6262.120996496496u,0 6262.121996496497u,1.5 6265.053616616617u,1.5 6265.054616616617u,0 6266.031156656657u,0 6266.032156656657u,1.5 6267.0086966966965u,1.5 6267.009696696697u,0 6268.963776776777u,0 6268.964776776777u,1.5 6269.941316816817u,1.5 6269.942316816817u,0 6270.918856856857u,0 6270.919856856857u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6273.851476976977u,0 6273.852476976977u,1.5 6274.829017017017u,1.5 6274.830017017017u,0 6275.806557057057u,0 6275.807557057057u,1.5 6276.784097097097u,1.5 6276.785097097098u,0 6277.761637137137u,0 6277.762637137137u,1.5 6279.716717217217u,1.5 6279.717717217217u,0 6282.649337337337u,0 6282.650337337337u,1.5 6283.626877377377u,1.5 6283.627877377377u,0 6284.604417417418u,0 6284.605417417418u,1.5 6287.537037537537u,1.5 6287.538037537537u,0 6288.514577577577u,0 6288.5155775775775u,1.5 6296.3348978978975u,1.5 6296.335897897898u,0 6298.289977977978u,0 6298.290977977978u,1.5 6300.245058058058u,1.5 6300.246058058058u,0 6304.155218218218u,0 6304.156218218218u,1.5 6305.132758258259u,1.5 6305.133758258259u,0 6309.042918418419u,0 6309.043918418419u,1.5 6310.020458458459u,1.5 6310.021458458459u,0 6313.930618618619u,0 6313.931618618619u,1.5 6314.908158658659u,1.5 6314.909158658659u,0 6315.885698698698u,0 6315.886698698699u,1.5 6317.840778778779u,1.5 6317.841778778779u,0 6318.818318818819u,0 6318.819318818819u,1.5 6319.795858858859u,1.5 6319.796858858859u,0 6320.773398898898u,0 6320.774398898899u,1.5 6321.750938938939u,1.5 6321.751938938939u,0 6326.638639139139u,0 6326.639639139139u,1.5 6329.57125925926u,1.5 6329.57225925926u,0 6330.548799299299u,0 6330.5497992993u,1.5 6331.526339339339u,1.5 6331.527339339339u,0 6337.391579579579u,0 6337.392579579579u,1.5 6339.34665965966u,1.5 6339.34765965966u,0 6340.324199699699u,0 6340.3251996997u,1.5 6342.27927977978u,1.5 6342.28027977978u,0 6343.25681981982u,0 6343.25781981982u,1.5 6344.23435985986u,1.5 6344.23535985986u,0 6350.0996001001u,0 6350.100600100101u,1.5 6351.07714014014u,1.5 6351.07814014014u,0 6352.05468018018u,0 6352.05568018018u,1.5 6354.009760260261u,1.5 6354.010760260261u,0 6354.9873003003u,0 6354.988300300301u,1.5 6355.96484034034u,1.5 6355.96584034034u,0 6356.94238038038u,0 6356.94338038038u,1.5 6358.897460460461u,1.5 6358.898460460461u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6363.785160660661u,0 6363.786160660661u,1.5 6370.627940940941u,1.5 6370.628940940941u,0 6371.605480980981u,0 6371.606480980981u,1.5 6372.583021021021u,1.5 6372.584021021021u,0 6379.425801301301u,0 6379.426801301302u,1.5 6386.268581581581u,1.5 6386.269581581581u,0 6388.223661661662u,0 6388.224661661662u,1.5 6389.201201701701u,1.5 6389.202201701702u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6397.021522022022u,0 6397.022522022022u,1.5 6397.999062062062u,1.5 6398.000062062062u,0 6398.976602102102u,0 6398.9776021021025u,1.5 6400.931682182182u,1.5 6400.932682182182u,0 6401.909222222222u,0 6401.910222222222u,1.5 6404.841842342342u,1.5 6404.842842342342u,0 6406.7969224224225u,0 6406.797922422423u,1.5 6407.774462462463u,1.5 6407.775462462463u,0 6410.707082582582u,0 6410.708082582582u,1.5 6411.684622622623u,1.5 6411.685622622623u,0 6414.617242742742u,0 6414.618242742742u,1.5 6416.572322822823u,1.5 6416.573322822823u,0 6417.549862862863u,0 6417.550862862863u,1.5 6420.482482982983u,1.5 6420.483482982983u,0 6421.460023023023u,0 6421.461023023023u,1.5 6422.437563063063u,1.5 6422.438563063063u,0 6426.347723223223u,0 6426.348723223223u,1.5 6427.325263263264u,1.5 6427.326263263264u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6437.100663663664u,0 6437.101663663664u,1.5 6445.898524024024u,1.5 6445.899524024024u,0 6448.831144144144u,0 6448.832144144144u,1.5 6449.808684184184u,1.5 6449.809684184184u,0 6451.763764264265u,0 6451.764764264265u,1.5 6452.741304304304u,1.5 6452.7423043043045u,0 6454.696384384384u,0 6454.697384384384u,1.5 6456.651464464465u,1.5 6456.652464464465u,0 6463.494244744744u,0 6463.495244744744u,1.5 6464.471784784785u,1.5 6464.472784784785u,0 6465.4493248248245u,0 6465.450324824825u,1.5 6466.426864864865u,1.5 6466.427864864865u,0 6468.381944944945u,0 6468.382944944945u,1.5 6469.359484984985u,1.5 6469.360484984985u,0 6471.314565065065u,0 6471.315565065065u,1.5 6472.292105105105u,1.5 6472.2931051051055u,0 6474.247185185185u,0 6474.248185185185u,1.5 6476.202265265266u,1.5 6476.203265265266u,0 6477.179805305305u,0 6477.1808053053055u,1.5 6484.022585585586u,1.5 6484.023585585586u,0 6485.0001256256255u,0 6485.001125625626u,1.5 6488.910285785786u,1.5 6488.911285785786u,0 6490.865365865866u,0 6490.866365865866u,1.5 6496.730606106106u,1.5 6496.7316061061065u,0 6497.708146146146u,0 6497.709146146146u,1.5 6500.640766266267u,1.5 6500.641766266267u,0 6501.618306306306u,0 6501.6193063063065u,1.5 6511.393706706706u,1.5 6511.3947067067065u,0 6512.371246746747u,0 6512.372246746747u,1.5 6513.348786786787u,1.5 6513.349786786787u,0 6514.3263268268265u,0 6514.327326826827u,1.5 6517.258946946947u,1.5 6517.259946946947u,0 6518.236486986987u,0 6518.237486986987u,1.5 6520.191567067067u,1.5 6520.192567067067u,0 6521.169107107107u,0 6521.1701071071075u,1.5 6525.079267267268u,1.5 6525.080267267268u,0 6527.034347347347u,0 6527.035347347347u,1.5 6528.9894274274275u,1.5 6528.990427427428u,0 6532.899587587588u,0 6532.900587587588u,1.5 6533.8771276276275u,1.5 6533.878127627628u,0 6535.832207707707u,0 6535.8332077077075u,1.5 6536.809747747748u,1.5 6536.810747747748u,0 6543.6525280280275u,0 6543.653528028028u,1.5 6544.630068068068u,1.5 6544.631068068068u,0 6549.517768268269u,0 6549.518768268269u,1.5 6551.472848348348u,1.5 6551.473848348348u,0 6553.4279284284285u,0 6553.428928428429u,1.5 6562.225788788789u,1.5 6562.226788788789u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6565.158408908908u,0 6565.1594089089085u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6568.0910290290285u,0 6568.092029029029u,1.5 6569.068569069069u,1.5 6569.069569069069u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.001189189189u,1.5 6572.002189189189u,0 6574.933809309309u,0 6574.9348093093095u,1.5 6575.911349349349u,1.5 6575.912349349349u,0 6577.866429429429u,0 6577.86742942943u,1.5 6586.66428978979u,1.5 6586.66528978979u,0 6587.6418298298295u,0 6587.64282982983u,1.5 6588.61936986987u,1.5 6588.62036986987u,0 6590.57444994995u,0 6590.57544994995u,1.5 6592.5295300300295u,1.5 6592.53053003003u,0 6596.43969019019u,0 6596.44069019019u,1.5 6597.4172302302295u,1.5 6597.41823023023u,0 6598.394770270271u,0 6598.395770270271u,1.5 6600.34985035035u,1.5 6600.35085035035u,0 6601.32739039039u,0 6601.32839039039u,1.5 6602.30493043043u,1.5 6602.305930430431u,0 6603.282470470471u,0 6603.283470470471u,1.5 6604.26001051051u,1.5 6604.2610105105105u,0 6606.215090590591u,0 6606.216090590591u,1.5 6607.19263063063u,1.5 6607.193630630631u,0 6612.0803308308305u,0 6612.081330830831u,1.5 6613.057870870871u,1.5 6613.058870870871u,0 6614.03541091091u,0 6614.0364109109105u,1.5 6615.012950950951u,1.5 6615.013950950951u,0 6615.990490990991u,0 6615.991490990991u,1.5 6617.945571071071u,1.5 6617.946571071071u,0 6619.900651151151u,0 6619.901651151151u,1.5 6621.8557312312305u,1.5 6621.856731231231u,0 6623.810811311311u,0 6623.811811311311u,1.5 6624.788351351351u,1.5 6624.789351351351u,0 6626.743431431431u,0 6626.744431431432u,1.5 6627.720971471472u,1.5 6627.721971471472u,0 6629.676051551551u,0 6629.677051551551u,1.5 6631.631131631631u,1.5 6631.632131631632u,0 6632.608671671672u,0 6632.609671671672u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6637.496371871872u,1.5 6637.497371871872u,0 6638.473911911911u,0 6638.4749119119115u,1.5 6639.451451951952u,1.5 6639.452451951952u,0 6643.361612112112u,0 6643.362612112112u,1.5 6645.316692192192u,1.5 6645.317692192192u,0 6646.2942322322315u,0 6646.295232232232u,1.5 6649.226852352352u,1.5 6649.227852352352u,0 6650.204392392392u,0 6650.205392392392u,1.5 6651.181932432432u,1.5 6651.182932432433u,0 6654.114552552552u,0 6654.115552552552u,1.5 6655.092092592593u,1.5 6655.093092592593u,0 6657.047172672673u,0 6657.048172672673u,1.5 6659.002252752753u,1.5 6659.003252752753u,0 6659.979792792793u,0 6659.980792792793u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6664.867492992993u,0 6664.868492992993u,1.5 6666.822573073073u,1.5 6666.823573073073u,0 6668.777653153153u,0 6668.778653153153u,1.5 6672.687813313313u,1.5 6672.688813313313u,0 6673.665353353353u,0 6673.666353353353u,1.5 6674.642893393393u,1.5 6674.643893393393u,0 6676.597973473474u,0 6676.598973473474u,1.5 6677.575513513513u,1.5 6677.576513513513u,0 6678.553053553553u,0 6678.554053553553u,1.5 6679.530593593594u,1.5 6679.531593593594u,0 6680.508133633633u,0 6680.509133633634u,1.5 6684.418293793794u,1.5 6684.419293793794u,0 6691.261074074074u,0 6691.262074074074u,1.5 6693.216154154154u,1.5 6693.217154154154u,0 6694.193694194194u,0 6694.194694194194u,1.5 6698.103854354354u,1.5 6698.104854354354u,0 6702.991554554554u,0 6702.992554554554u,1.5 6704.946634634634u,1.5 6704.947634634635u,0 6706.901714714714u,0 6706.902714714714u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6708.856794794795u,0 6708.857794794795u,1.5 6709.834334834834u,1.5 6709.835334834835u,0 6711.789414914914u,0 6711.790414914914u,1.5 6712.766954954955u,1.5 6712.767954954955u,0 6713.744494994995u,0 6713.745494994995u,1.5 6715.699575075075u,1.5 6715.700575075075u,0 6716.677115115115u,0 6716.678115115115u,1.5 6718.632195195195u,1.5 6718.633195195195u,0 6719.609735235234u,0 6719.610735235235u,1.5 6720.587275275276u,1.5 6720.588275275276u,0 6723.519895395395u,0 6723.520895395395u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6727.430055555555u,0 6727.431055555555u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6733.295295795796u,0 6733.296295795796u,1.5 6734.272835835835u,1.5 6734.273835835836u,0 6735.250375875876u,0 6735.251375875876u,1.5 6736.227915915916u,1.5 6736.228915915916u,0 6737.205455955956u,0 6737.206455955956u,1.5 6741.115616116116u,1.5 6741.116616116116u,0 6742.093156156156u,0 6742.094156156156u,1.5 6743.070696196196u,1.5 6743.071696196196u,0 6744.048236236235u,0 6744.049236236236u,1.5 6745.025776276277u,1.5 6745.026776276277u,0 6746.003316316316u,0 6746.004316316316u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6753.823636636636u,1.5 6753.824636636637u,0 6754.801176676677u,0 6754.802176676677u,1.5 6761.6439569569575u,1.5 6761.644956956958u,0 6766.5316571571575u,0 6766.532657157158u,1.5 6768.486737237236u,1.5 6768.487737237237u,0 6769.464277277278u,0 6769.465277277278u,1.5 6771.4193573573575u,1.5 6771.420357357358u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6775.329517517517u,0 6775.330517517517u,1.5 6776.3070575575575u,1.5 6776.308057557558u,0 6777.284597597598u,0 6777.285597597598u,1.5 6778.262137637637u,1.5 6778.263137637638u,0 6779.239677677678u,0 6779.240677677678u,1.5 6780.217217717717u,1.5 6780.218217717717u,0 6782.172297797798u,0 6782.173297797798u,1.5 6783.149837837837u,1.5 6783.150837837838u,0 6786.0824579579585u,0 6786.083457957959u,1.5 6787.059997997998u,1.5 6787.060997997998u,0 6788.037538038037u,0 6788.038538038038u,1.5 6791.947698198198u,1.5 6791.948698198198u,0 6794.880318318318u,0 6794.881318318318u,1.5 6795.8578583583585u,1.5 6795.858858358359u,0 6798.790478478479u,0 6798.791478478479u,1.5 6802.700638638638u,1.5 6802.7016386386385u,0 6803.678178678679u,0 6803.679178678679u,1.5 6805.633258758759u,1.5 6805.63425875876u,0 6808.565878878879u,0 6808.566878878879u,1.5 6810.520958958959u,1.5 6810.52195895896u,0 6811.498498998999u,0 6811.499498998999u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6814.431119119119u,0 6814.432119119119u,1.5 6815.4086591591595u,1.5 6815.40965915916u,0 6818.34127927928u,0 6818.34227927928u,1.5 6819.318819319319u,1.5 6819.319819319319u,0 6821.273899399399u,0 6821.274899399399u,1.5 6823.22897947948u,1.5 6823.22997947948u,0 6824.206519519519u,0 6824.207519519519u,1.5 6826.1615995996u,1.5 6826.1625995996u,0 6827.139139639639u,0 6827.1401396396395u,1.5 6828.11667967968u,1.5 6828.11767967968u,0 6831.0492997998u,0 6831.0502997998u,1.5 6832.026839839839u,1.5 6832.0278398398395u,0 6833.00437987988u,0 6833.00537987988u,1.5 6833.98191991992u,1.5 6833.98291991992u,0 6834.95945995996u,0 6834.960459959961u,1.5 6835.937u,1.5 6835.938u,0 6837.89208008008u,0 6837.89308008008u,1.5 6839.8471601601605u,1.5 6839.848160160161u,0 6841.802240240239u,0 6841.80324024024u,1.5 6842.779780280281u,1.5 6842.780780280281u,0 6844.7348603603605u,0 6844.735860360361u,1.5 6845.7124004004u,1.5 6845.7134004004u,0 6846.68994044044u,0 6846.6909404404405u,1.5 6848.64502052052u,1.5 6848.64602052052u,0 6849.6225605605605u,0 6849.623560560561u,1.5 6851.57764064064u,1.5 6851.5786406406405u,0 6854.510260760761u,0 6854.511260760762u,1.5 6856.46534084084u,1.5 6856.4663408408405u,0 6857.442880880881u,0 6857.443880880881u,1.5 6859.397960960961u,1.5 6859.398960960962u,0 6861.35304104104u,0 6861.354041041041u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6866.24074124124u,0 6866.241741241241u,1.5 6867.218281281282u,1.5 6867.219281281282u,0 6870.150901401401u,0 6870.151901401401u,1.5 6871.128441441441u,1.5 6871.1294414414415u,0 6872.105981481482u,0 6872.106981481482u,1.5 6876.016141641641u,1.5 6876.0171416416415u,0 6876.993681681682u,0 6876.994681681682u,1.5 6878.948761761762u,1.5 6878.949761761763u,0 6884.814002002002u,0 6884.815002002002u,1.5 6885.791542042041u,1.5 6885.7925420420415u,0 6886.769082082082u,0 6886.770082082082u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6893.611862362362u,0 6893.612862362363u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6900.454642642642u,0 6900.4556426426425u,1.5 6901.432182682683u,1.5 6901.433182682683u,0 6903.387262762763u,0 6903.388262762764u,1.5 6907.297422922923u,1.5 6907.298422922923u,0 6909.252503003003u,0 6909.253503003003u,1.5 6912.185123123123u,1.5 6912.186123123123u,0 6913.162663163163u,0 6913.163663163164u,1.5 6914.140203203203u,1.5 6914.141203203203u,0 6920.982983483484u,0 6920.983983483484u,1.5 6922.938063563563u,1.5 6922.939063563564u,0 6924.893143643643u,0 6924.8941436436435u,1.5 6926.848223723723u,1.5 6926.849223723723u,0 6927.825763763764u,0 6927.826763763765u,1.5 6932.713463963964u,1.5 6932.714463963965u,0 6933.691004004004u,0 6933.692004004004u,1.5 6934.668544044043u,1.5 6934.6695440440435u,0 6935.646084084084u,0 6935.647084084084u,1.5 6936.623624124124u,1.5 6936.624624124124u,0 6938.578704204204u,0 6938.579704204204u,1.5 6939.556244244243u,1.5 6939.5572442442435u,0 6942.488864364364u,0 6942.489864364365u,1.5 6943.466404404404u,1.5 6943.467404404404u,0 6945.421484484485u,0 6945.422484484485u,1.5 6946.399024524524u,1.5 6946.400024524524u,0 6950.309184684685u,0 6950.310184684685u,1.5 6954.219344844844u,1.5 6954.2203448448445u,0 6955.196884884885u,0 6955.197884884885u,1.5 6958.129505005005u,1.5 6958.130505005005u,0 6959.107045045044u,0 6959.1080450450445u,1.5 6962.039665165165u,1.5 6962.040665165166u,0 6963.017205205205u,0 6963.018205205205u,1.5 6963.994745245244u,1.5 6963.9957452452445u,0 6964.972285285286u,0 6964.973285285286u,1.5 6967.904905405405u,1.5 6967.905905405405u,0 6968.882445445445u,0 6968.883445445445u,1.5 6969.859985485486u,1.5 6969.860985485486u,0 6970.837525525525u,0 6970.838525525525u,1.5 6971.815065565565u,1.5 6971.816065565566u,0 6972.792605605606u,0 6972.793605605606u,1.5 6973.770145645645u,1.5 6973.771145645645u,0 6974.747685685686u,0 6974.748685685686u,1.5 6976.702765765766u,1.5 6976.703765765767u,0 6978.657845845845u,0 6978.6588458458455u,1.5 6980.612925925926u,1.5 6980.613925925926u,0 6981.590465965966u,0 6981.591465965967u,1.5 6982.568006006006u,1.5 6982.569006006006u,0 6986.478166166166u,0 6986.479166166167u,1.5 6987.455706206206u,1.5 6987.456706206206u,0 6988.433246246245u,0 6988.4342462462455u,1.5 6990.388326326326u,1.5 6990.389326326326u,0 6991.365866366366u,0 6991.366866366367u,1.5 6992.343406406406u,1.5 6992.344406406406u,0 6994.298486486487u,0 6994.299486486487u,1.5 6995.276026526526u,1.5 6995.277026526526u,0
vbb12 bb12 0 pwl 0,1.5  3.90966016016016u,1.5 3.9106601601601603u,0 4.8872002002002u,0 4.8882002002002u,1.5 10.75244044044044u,1.5 10.753440440440441u,0 11.72998048048048u,0 11.730980480480481u,1.5 12.70752052052052u,1.5 12.708520520520521u,0 13.68506056056056u,0 13.686060560560561u,1.5 17.59522072072072u,1.5 17.59622072072072u,0 18.572760760760765u,0 18.573760760760763u,1.5 25.415541041041042u,1.5 25.41654104104104u,0 26.393081081081085u,0 26.394081081081083u,1.5 27.370621121121122u,1.5 27.37162112112112u,0 28.348161161161162u,0 28.34916116116116u,1.5 30.303241241241246u,1.5 30.304241241241243u,0 31.280781281281282u,0 31.28178128128128u,1.5 33.23586136136136u,1.5 33.23686136136136u,0 35.19094144144144u,0 35.19194144144144u,1.5 36.16848148148148u,1.5 36.16948148148148u,0 37.146021521521526u,0 37.14702152152153u,1.5 38.12356156156156u,1.5 38.12456156156156u,0 40.07864164164164u,0 40.07964164164164u,1.5 41.05618168168168u,1.5 41.05718168168168u,0 58.6519024024024u,0 58.652902402402404u,1.5 59.62944244244244u,1.5 59.630442442442444u,0 63.539602602602606u,0 63.54060260260261u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 85.04548348348348u,1.5 85.04648348348348u,0 86.02302352352352u,0 86.02402352352352u,1.5 87.00056356356356u,1.5 87.00156356356356u,0 90.91072372372372u,0 90.91172372372372u,1.5 91.88826376376376u,1.5 91.88926376376376u,0 104.59628428428428u,0 104.59728428428429u,1.5 106.55136436436436u,1.5 106.55236436436437u,0 107.5289044044044u,0 107.5299044044044u,1.5 109.48398448448448u,1.5 109.48498448448449u,0 110.46152452452452u,0 110.46252452452453u,1.5 116.32676476476476u,1.5 116.32776476476477u,0 117.3043048048048u,0 117.3053048048048u,1.5 123.16954504504503u,1.5 123.17054504504503u,0 124.14708508508508u,0 124.14808508508509u,1.5 125.12462512512512u,1.5 125.12562512512513u,0 135.8775655655656u,0 135.87856556556557u,1.5 136.85510560560562u,1.5 136.8561056056056u,0 137.83264564564567u,0 137.83364564564565u,1.5 150.54066616616618u,1.5 150.54166616616615u,0 152.49574624624626u,0 152.49674624624623u,1.5 153.4732862862863u,1.5 153.4742862862863u,0 158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 164.22622672672674u,0 164.2272267267267u,1.5 174.97916716716716u,1.5 174.98016716716714u,0 184.7545675675676u,0 184.75556756756757u,1.5 185.73210760760762u,1.5 185.7331076076076u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 188.66472772772775u,0 188.66572772772773u,1.5 195.50750800800802u,1.5 195.508508008008u,0 197.4625880880881u,0 197.46358808808807u,1.5 198.44012812812815u,1.5 198.44112812812813u,0 207.2379884884885u,0 207.23898848848847u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 210.17060860860863u,0 210.1716086086086u,1.5 218.96846896896898u,1.5 218.96946896896895u,0 219.94600900900903u,0 219.947009009009u,1.5 220.92354904904906u,1.5 220.92454904904903u,0 229.72140940940943u,0 229.7224094094094u,1.5 230.69894944944946u,1.5 230.69994944944943u,0 231.6764894894895u,0 231.6774894894895u,1.5 237.54172972972972u,1.5 237.5427297297297u,0 238.51926976976978u,0 238.52026976976975u,1.5 239.4968098098098u,1.5 239.49780980980978u,0 240.47434984984986u,0 240.47534984984983u,1.5 241.4518898898899u,1.5 241.4528898898899u,0 242.42942992992997u,0 242.43042992992994u,1.5 243.40696996996996u,1.5 243.40796996996994u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 259.04761061061066u,1.5 259.04861061061064u,0 260.02515065065063u,0 260.0261506506506u,1.5 261.00269069069066u,1.5 261.00369069069063u,0 261.98023073073074u,0 261.9812307307307u,1.5 262.95777077077076u,1.5 262.95877077077074u,0 270.77809109109114u,0 270.7790910910911u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 272.73317117117114u,0 272.7341711711711u,1.5 279.57595145145143u,1.5 279.5769514514514u,0 280.5534914914915u,0 280.5544914914915u,1.5 281.53103153153154u,1.5 281.5320315315315u,0 282.50857157157157u,0 282.50957157157154u,1.5 283.48611161161165u,1.5 283.4871116116116u,0 289.35135185185186u,0 289.35235185185184u,1.5 290.32889189189194u,1.5 290.3298918918919u,0 294.23905205205205u,0 294.240052052052u,1.5 302.0593723723724u,1.5 302.0603723723724u,0 304.0144524524524u,0 304.0154524524524u,1.5 305.9695325325325u,1.5 305.9705325325325u,0 306.9470725725726u,0 306.9480725725726u,1.5 307.92461261261263u,1.5 307.9256126126126u,0 313.78985285285285u,0 313.7908528528528u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 315.74493293293295u,0 315.74593293293293u,1.5 317.700013013013u,1.5 317.701013013013u,0 318.67755305305303u,0 318.678553053053u,1.5 323.5652532532532u,1.5 323.5662532532532u,0 324.5427932932933u,0 324.5437932932933u,1.5 326.4978733733734u,1.5 326.4988733733734u,0 328.45295345345346u,0 328.45395345345344u,1.5 329.4304934934935u,1.5 329.43149349349346u,0 335.2957337337337u,0 335.2967337337337u,1.5 336.2732737737738u,1.5 336.27427377377376u,0 337.2508138138138u,0 337.2518138138138u,1.5 338.2283538538539u,1.5 338.22935385385387u,0 340.18343393393394u,0 340.1844339339339u,1.5 349.9588343343343u,1.5 349.9598343343343u,0 350.9363743743744u,0 350.9373743743744u,1.5 351.9139144144144u,1.5 351.9149144144144u,0 352.8914544544545u,0 352.8924544544545u,1.5 353.8689944944945u,1.5 353.86999449449445u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 374.39733533533536u,1.5 374.39833533533533u,0 375.3748753753754u,0 375.37587537537536u,1.5 378.3074954954955u,1.5 378.3084954954955u,0 380.26257557557557u,0 380.26357557557554u,1.5 381.2401156156156u,1.5 381.24111561561557u,0 389.06043593593597u,0 389.06143593593595u,1.5 390.037975975976u,1.5 390.038975975976u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 395.90321621621626u,0 395.90421621621624u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 405.67861661661664u,1.5 405.6796166166166u,0 406.65615665665666u,0 406.65715665665664u,1.5 408.61123673673677u,1.5 408.61223673673675u,0 409.5887767767768u,0 409.5897767767768u,1.5 410.5663168168168u,1.5 410.5673168168168u,0 411.54385685685685u,0 411.5448568568568u,1.5 412.5213968968969u,1.5 412.52239689689685u,0 414.476476976977u,0 414.47747697697696u,1.5 415.45401701701707u,1.5 415.45501701701704u,0 432.07219769769773u,0 432.0731976976977u,1.5 433.04973773773776u,1.5 433.05073773773773u,0 434.0272777777778u,0 434.02827777777776u,1.5 435.00481781781787u,1.5 435.00581781781784u,0 435.98235785785783u,0 435.9833578578578u,1.5 437.93743793793794u,1.5 437.9384379379379u,0 438.91497797797797u,0 438.91597797797795u,1.5 455.53315865865864u,1.5 455.5341586586586u,0 456.5106986986987u,0 456.5116986986987u,1.5 462.37593893893893u,1.5 462.3769389389389u,0 463.353478978979u,0 463.354478978979u,1.5 466.28609909909915u,1.5 466.2870990990991u,0 468.2411791791792u,0 468.2421791791792u,1.5 470.19625925925925u,1.5 470.1972592592592u,0 471.17379929929933u,0 471.1747992992993u,1.5 472.15133933933936u,1.5 472.15233933933933u,0 474.1064194194194u,0 474.1074194194194u,1.5 475.08395945945944u,1.5 475.0849594594594u,0 476.0614994994995u,0 476.0624994994995u,1.5 478.0165795795796u,1.5 478.0175795795796u,0 486.8144399399399u,0 486.8154399399399u,1.5 487.79197997998u,1.5 487.79297997998u,0 488.7695200200201u,0 488.77052002002006u,1.5 489.7470600600601u,1.5 489.7480600600601u,0 496.58984034034034u,0 496.5908403403403u,1.5 497.56738038038037u,1.5 497.56838038038035u,0 503.4326206206207u,0 503.4336206206207u,1.5 504.41016066066067u,1.5 504.41116066066064u,0 509.2978608608609u,0 509.2988608608609u,1.5 510.2754009009009u,1.5 510.27640090090085u,0 518.0957212212213u,0 518.0967212212213u,1.5 519.0732612612613u,1.5 519.0742612612613u,0 521.0283413413413u,0 521.0293413413413u,1.5 522.0058813813813u,1.5 522.0068813813813u,0 525.9160415415415u,0 525.9170415415415u,1.5 526.8935815815815u,1.5 526.8945815815815u,0 528.8486616616617u,0 528.8496616616617u,1.5 530.8037417417418u,1.5 530.8047417417417u,0 531.7812817817818u,0 531.7822817817818u,1.5 533.7363618618618u,1.5 533.7373618618618u,0 534.7139019019019u,0 534.7149019019018u,1.5 540.5791421421421u,1.5 540.5801421421421u,0 541.5566821821823u,0 541.5576821821822u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 561.107482982983u,0 561.108482982983u,1.5 563.0625630630631u,1.5 563.063563063063u,0 564.0401031031031u,0 564.0411031031031u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 568.9278033033033u,0 568.9288033033033u,1.5 569.9053433433434u,1.5 569.9063433433433u,0 584.5684439439439u,0 584.5694439439438u,1.5 585.545983983984u,1.5 585.546983983984u,0 587.501064064064u,0 587.502064064064u,1.5 589.4561441441441u,1.5 589.4571441441441u,0 590.4336841841842u,0 590.4346841841842u,1.5 592.3887642642643u,1.5 592.3897642642643u,0 593.3663043043043u,0 593.3673043043043u,1.5 596.2989244244244u,1.5 596.2999244244244u,0 597.2764644644644u,0 597.2774644644644u,1.5 602.1641646646647u,1.5 602.1651646646646u,0 603.1417047047047u,0 603.1427047047047u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 606.0743248248249u,0 606.0753248248249u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 620.7374254254254u,0 620.7384254254254u,1.5 621.7149654654654u,1.5 621.7159654654654u,0 623.6700455455456u,0 623.6710455455456u,1.5 637.355606106106u,1.5 637.356606106106u,0 649.0860865865866u,0 649.0870865865866u,1.5 660.816567067067u,1.5 660.817567067067u,0 661.7941071071072u,0 661.7951071071071u,1.5 662.7716471471472u,1.5 662.7726471471472u,0 663.7491871871872u,0 663.7501871871872u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 672.5470475475475u,0 672.5480475475475u,1.5 674.5021276276276u,1.5 674.5031276276276u,0 675.4796676676676u,0 675.4806676676676u,1.5 685.255068068068u,1.5 685.256068068068u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 696.0080085085085u,0 696.0090085085085u,1.5 696.9855485485485u,1.5 696.9865485485485u,0 697.9630885885886u,0 697.9640885885885u,1.5 707.7384889889889u,1.5 707.7394889889889u,0 708.716029029029u,0 708.7170290290289u,1.5 709.693569069069u,1.5 709.694569069069u,0 716.5363493493494u,0 716.5373493493494u,1.5 717.5138893893894u,1.5 717.5148893893894u,0 718.4914294294294u,0 718.4924294294294u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 729.24436986987u,1.5 729.2453698698699u,0 730.22190990991u,0 730.22290990991u,1.5 731.19944994995u,1.5 731.20044994995u,0 739.0197702702703u,0 739.0207702702703u,1.5 740.9748503503504u,1.5 740.9758503503504u,0 741.9523903903904u,0 741.9533903903904u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 761.5031911911911u,0 761.5041911911911u,1.5 762.4807312312312u,1.5 762.4817312312312u,0 763.4582712712713u,0 763.4592712712713u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 771.2785915915915u,0 771.2795915915915u,1.5 772.2561316316315u,1.5 772.2571316316315u,0 781.053991991992u,0 781.054991991992u,1.5 782.031532032032u,1.5 782.032532032032u,0 783.0090720720721u,0 783.010072072072u,1.5 790.8293923923924u,1.5 790.8303923923924u,0 792.7844724724725u,0 792.7854724724725u,1.5 793.7620125125126u,1.5 793.7630125125125u,0 803.5374129129129u,0 803.5384129129129u,1.5 814.2903533533533u,1.5 814.2913533533533u,0 815.2678933933934u,0 815.2688933933933u,1.5 816.2454334334335u,1.5 816.2464334334335u,0 825.0432937937937u,0 825.0442937937937u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 841.6614744744745u,1.5 841.6624744744745u,0 848.5042547547547u,0 848.5052547547547u,1.5 849.4817947947948u,1.5 849.4827947947948u,0 851.4368748748749u,0 851.4378748748749u,1.5 854.3694949949951u,1.5 854.370494994995u,0 855.3470350350351u,0 855.3480350350351u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 868.0550555555556u,0 868.0560555555555u,1.5 869.0325955955957u,1.5 869.0335955955957u,0 878.8079959959961u,0 878.808995995996u,1.5 894.4486366366367u,1.5 894.4496366366367u,0 896.4037167167166u,0 896.4047167167166u,1.5 897.3812567567567u,1.5 897.3822567567566u,0 908.1341971971972u,0 908.1351971971972u,1.5 909.1117372372372u,1.5 909.1127372372372u,0 911.0668173173173u,0 911.0678173173172u,1.5 912.0443573573574u,1.5 912.0453573573574u,0 913.0218973973974u,0 913.0228973973974u,1.5 913.9994374374375u,1.5 914.0004374374374u,0 914.9769774774775u,0 914.9779774774775u,1.5 916.9320575575576u,1.5 916.9330575575576u,0 917.9095975975977u,0 917.9105975975976u,1.5 927.684997997998u,1.5 927.685997997998u,0 928.6625380380381u,0 928.663538038038u,1.5 932.5726981981983u,1.5 932.5736981981983u,0 933.5502382382382u,0 933.5512382382382u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 938.4379384384384u,0 938.4389384384384u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 959.9438193193192u,0 959.9448193193192u,1.5 960.9213593593594u,1.5 960.9223593593593u,0 964.8315195195195u,0 964.8325195195195u,1.5 966.7865995995996u,1.5 966.7875995995996u,0 967.7641396396397u,0 967.7651396396396u,1.5 968.7416796796797u,1.5 968.7426796796797u,0 970.6967597597597u,0 970.6977597597597u,1.5 972.6518398398398u,1.5 972.6528398398398u,0 973.6293798798798u,0 973.6303798798798u,1.5 974.60691991992u,1.5 974.6079199199199u,0 975.58445995996u,0 975.58545995996u,1.5 977.5395400400402u,1.5 977.5405400400401u,0 978.5170800800801u,0 978.51808008008u,1.5 981.4497002002003u,1.5 981.4507002002002u,0 982.4272402402403u,0 982.4282402402403u,1.5 983.4047802802802u,1.5 983.4057802802802u,0 984.3823203203203u,0 984.3833203203203u,1.5 989.2700205205206u,1.5 989.2710205205206u,0 990.2475605605605u,0 990.2485605605605u,1.5 991.2251006006006u,1.5 991.2261006006006u,0 992.2026406406408u,0 992.2036406406407u,1.5 994.1577207207208u,1.5 994.1587207207208u,0 995.1352607607607u,0 995.1362607607607u,1.5 999.045420920921u,1.5 999.0464209209209u,0 1000.0229609609609u,0 1000.0239609609608u,1.5 1001.9780410410411u,1.5 1001.9790410410411u,0 1002.955581081081u,0 1002.956581081081u,1.5 1004.9106611611611u,1.5 1004.9116611611611u,0 1005.8882012012012u,0 1005.8892012012012u,1.5 1013.7085215215216u,1.5 1013.7095215215215u,0 1014.6860615615615u,0 1014.6870615615614u,1.5 1016.6411416416418u,1.5 1016.6421416416417u,0 1017.6186816816817u,0 1017.6196816816816u,1.5 1021.5288418418419u,1.5 1021.5298418418419u,0 1022.5063818818818u,0 1022.5073818818818u,1.5 1026.416542042042u,1.5 1026.4175420420422u,0 1027.394082082082u,0 1027.3950820820821u,1.5 1028.371622122122u,1.5 1028.3726221221223u,0 1029.349162162162u,0 1029.3501621621622u,1.5 1030.3267022022021u,1.5 1030.3277022022023u,0 1031.3042422422423u,0 1031.3052422422425u,1.5 1032.2817822822822u,1.5 1032.2827822822824u,0 1033.2593223223223u,0 1033.2603223223225u,1.5 1034.2368623623622u,1.5 1034.2378623623624u,0 1057.6978233233233u,0 1057.6988233233235u,1.5 1058.6753633633632u,1.5 1058.6763633633634u,0 1061.6079834834834u,0 1061.6089834834836u,1.5 1062.5855235235235u,1.5 1062.5865235235237u,0 1065.5181436436435u,0 1065.5191436436437u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1070.4058438438437u,1.5 1070.406843843844u,0 1071.3833838838837u,0 1071.3843838838839u,1.5 1086.0464844844844u,1.5 1086.0474844844846u,0 1087.0240245245245u,0 1087.0250245245247u,1.5 1088.9791046046046u,1.5 1088.9801046046048u,0 1089.9566446446445u,0 1089.9576446446447u,1.5 1091.9117247247245u,1.5 1091.9127247247247u,0 1092.8892647647647u,0 1092.8902647647649u,1.5 1093.8668048048046u,1.5 1093.8678048048048u,0 1102.6646651651652u,0 1102.6656651651654u,1.5 1103.642205205205u,1.5 1103.6432052052053u,0 1104.6197452452452u,0 1104.6207452452454u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1107.5523653653654u,0 1107.5533653653656u,1.5 1108.5299054054053u,1.5 1108.5309054054055u,0 1109.5074454454455u,0 1109.5084454454457u,1.5 1120.2603858858856u,1.5 1120.2613858858858u,0 1121.2379259259258u,0 1121.238925925926u,1.5 1122.215465965966u,1.5 1122.216465965966u,0 1124.170546046046u,0 1124.1715460460462u,1.5 1125.1480860860859u,1.5 1125.149086086086u,0 1134.9234864864864u,0 1134.9244864864866u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1148.609047047047u,1.5 1148.6100470470471u,0 1150.564127127127u,0 1150.5651271271272u,1.5 1151.5416671671671u,1.5 1151.5426671671673u,0 1152.519207207207u,0 1152.5202072072072u,1.5 1153.4967472472472u,1.5 1153.4977472472474u,0 1154.474287287287u,0 1154.4752872872873u,1.5 1155.4518273273272u,1.5 1155.4528273273274u,0 1161.3170675675676u,0 1161.3180675675678u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1163.2721476476477u,0 1163.2731476476479u,1.5 1164.2496876876876u,1.5 1164.2506876876878u,0 1165.2272277277275u,0 1165.2282277277277u,1.5 1172.0700080080078u,1.5 1172.071008008008u,0 1173.047548048048u,0 1173.0485480480481u,1.5 1175.002628128128u,1.5 1175.0036281281282u,0 1177.9352482482482u,0 1177.9362482482484u,1.5 1178.912788288288u,1.5 1178.9137882882883u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1197.486049049049u,1.5 1197.4870490490491u,0 1199.441129129129u,0 1199.4421291291292u,1.5 1200.418669169169u,1.5 1200.4196691691693u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1208.2389894894895u,1.5 1208.2399894894897u,0 1210.1940695695696u,0 1210.1950695695698u,1.5 1217.0368498498497u,1.5 1217.0378498498499u,0 1218.0143898898898u,0 1218.01538988989u,1.5 1218.9919299299297u,1.5 1218.99292992993u,0 1219.9694699699699u,0 1219.97046996997u,1.5 1220.9470100100098u,1.5 1220.94801001001u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1231.6999504504504u,0 1231.7009504504506u,1.5 1241.4753508508506u,1.5 1241.4763508508508u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1254.1833713713713u,0 1254.1843713713715u,1.5 1260.0486116116115u,1.5 1260.0496116116117u,0 1261.0261516516516u,0 1261.0271516516518u,1.5 1262.0036916916918u,1.5 1262.004691691692u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1269.8240120120117u,1.5 1269.825012012012u,0 1270.8015520520519u,0 1270.802552052052u,1.5 1271.779092092092u,1.5 1271.7800920920922u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1280.5769524524524u,1.5 1280.5779524524526u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1291.3298928928928u,1.5 1291.330892892893u,0 1292.3074329329327u,0 1292.3084329329329u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1303.0603733733733u,1.5 1303.0613733733735u,0 1305.0154534534533u,0 1305.0164534534536u,1.5 1305.9929934934935u,1.5 1305.9939934934937u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1315.7683938938937u,1.5 1315.769393893894u,0 1316.7459339339337u,0 1316.7469339339339u,1.5 1327.4988743743743u,1.5 1327.4998743743745u,0 1329.4539544544543u,0 1329.4549544544545u,1.5 1330.4314944944945u,1.5 1330.4324944944947u,0 1338.251814814815u,0 1338.252814814815u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1342.1619749749748u,0 1342.162974974975u,1.5 1348.0272152152152u,1.5 1348.0282152152154u,0 1349.004755255255u,0 1349.0057552552553u,1.5 1350.9598353353351u,1.5 1350.9608353353353u,0 1352.9149154154154u,0 1352.9159154154156u,1.5 1353.8924554554553u,1.5 1353.8934554554555u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1367.578016016016u,1.5 1367.579016016016u,0 1368.5555560560558u,0 1368.556556056056u,1.5 1376.3758763763763u,1.5 1376.3768763763765u,0 1377.3534164164164u,0 1377.3544164164166u,1.5 1378.3309564564563u,1.5 1378.3319564564565u,0 1379.3084964964964u,0 1379.3094964964966u,1.5 1380.2860365365364u,1.5 1380.2870365365366u,0 1384.1961966966967u,0 1384.197196696697u,1.5 1385.1737367367366u,1.5 1385.1747367367368u,0 1392.016517017017u,0 1392.017517017017u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1400.8143773773772u,1.5 1400.8153773773774u,0 1401.7919174174174u,0 1401.7929174174176u,1.5 1408.6346976976977u,1.5 1408.6356976976979u,0 1409.6122377377376u,0 1409.6132377377378u,1.5 1411.5673178178179u,1.5 1411.568317817818u,0 1414.4999379379378u,0 1414.500937937938u,1.5 1415.4774779779777u,1.5 1415.478477977978u,0 1431.1181186186186u,0 1431.1191186186188u,1.5 1432.0956586586585u,1.5 1432.0966586586587u,0 1433.0731986986987u,0 1433.0741986986989u,1.5 1434.0507387387386u,1.5 1434.0517387387388u,0 1436.0058188188189u,0 1436.006818818819u,1.5 1438.938438938939u,1.5 1438.9394389389392u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1464.35447997998u,1.5 1464.3554799799801u,0 1465.3320200200199u,0 1465.33302002002u,1.5 1467.2871001001u,1.5 1467.2881001001u,0 1468.26464014014u,0 1468.2656401401402u,1.5 1470.21972022022u,1.5 1470.2207202202203u,0 1471.19726026026u,0 1471.1982602602602u,1.5 1473.1523403403403u,1.5 1473.1533403403405u,0 1474.1298803803802u,0 1474.1308803803804u,1.5 1476.0849604604603u,1.5 1476.0859604604605u,0 1477.0625005005004u,0 1477.0635005005006u,1.5 1478.0400405405405u,1.5 1478.0410405405407u,0 1480.9726606606605u,0 1480.9736606606607u,1.5 1481.9502007007006u,1.5 1481.9512007007008u,0 1482.9277407407408u,0 1482.928740740741u,1.5 1483.9052807807807u,1.5 1483.906280780781u,0 1494.658221221221u,0 1494.6592212212213u,1.5 1495.635761261261u,1.5 1495.6367612612612u,0 1513.231481981982u,0 1513.2324819819821u,1.5 1514.209022022022u,1.5 1514.2100220220223u,0 1520.074262262262u,0 1520.0752622622622u,1.5 1521.0518023023021u,1.5 1521.0528023023023u,0 1522.0293423423423u,0 1522.0303423423425u,1.5 1523.0068823823822u,1.5 1523.0078823823824u,0 1524.9619624624622u,0 1524.9629624624624u,1.5 1525.9395025025024u,1.5 1525.9405025025026u,0 1526.9170425425425u,0 1526.9180425425427u,1.5 1527.8945825825824u,1.5 1527.8955825825826u,0 1530.8272027027026u,0 1530.8282027027028u,1.5 1531.8047427427427u,1.5 1531.805742742743u,0 1532.7822827827827u,0 1532.7832827827829u,1.5 1562.108483983984u,1.5 1562.109483983984u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1565.041104104104u,1.5 1565.0421041041043u,0 1566.996184184184u,0 1566.997184184184u,1.5 1567.973724224224u,1.5 1567.9747242242242u,0 1579.7042047047046u,0 1579.7052047047048u,1.5 1580.6817447447447u,1.5 1580.682744744745u,0 1581.6592847847846u,0 1581.6602847847848u,1.5 1582.6368248248248u,1.5 1582.637824824825u,0 1583.614364864865u,0 1583.6153648648651u,1.5 1584.5919049049048u,1.5 1584.592904904905u,0 1586.5469849849849u,0 1586.547984984985u,1.5 1587.524525025025u,1.5 1587.5255250250252u,0 1589.479605105105u,0 1589.4806051051053u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1603.1651656656657u,0 1603.1661656656659u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1607.0753258258258u,1.5 1607.076325825826u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1618.805806306306u,0 1618.8068063063063u,1.5 1619.7833463463462u,1.5 1619.7843463463464u,0 1621.7384264264263u,0 1621.7394264264265u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1650.0870875875873u,0 1650.0880875875876u,1.5 1651.0646276276275u,1.5 1651.0656276276277u,0 1652.0421676676676u,0 1652.0431676676678u,1.5 1662.795108108108u,1.5 1662.7961081081082u,0 1674.5255885885883u,0 1674.5265885885885u,1.5 1675.5031286286285u,1.5 1675.5041286286287u,0 1676.4806686686686u,0 1676.4816686686688u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1689.1886891891893u,0 1689.1896891891895u,1.5 1690.1662292292292u,1.5 1690.1672292292294u,0 1695.0539294294292u,0 1695.0549294294294u,1.5 1696.0314694694694u,1.5 1696.0324694694696u,0 1698.9640895895895u,0 1698.9650895895898u,1.5 1704.8293298298297u,1.5 1704.83032982983u,0 1705.8068698698698u,0 1705.80786986987u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1719.4924304304302u,0 1719.4934304304304u,1.5 1728.2902907907908u,1.5 1728.291290790791u,0 1729.2678308308307u,0 1729.268830830831u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1737.0881511511511u,0 1737.0891511511513u,1.5 1738.0656911911913u,1.5 1738.0666911911915u,0 1740.998311311311u,0 1740.9993113113112u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1752.7287917917918u,1.5 1752.729791791792u,0 1758.594032032032u,0 1758.5950320320321u,1.5 1759.571572072072u,1.5 1759.5725720720723u,0 1761.526652152152u,0 1761.5276521521523u,1.5 1767.3918923923923u,1.5 1767.3928923923925u,0 1768.3694324324322u,0 1768.3704324324324u,1.5 1771.3020525525524u,1.5 1771.3030525525526u,0 1781.0774529529529u,0 1781.078452952953u,1.5 1784.010073073073u,1.5 1784.0110730730732u,0 1784.987613113113u,0 1784.9886131131132u,1.5 1790.852853353353u,1.5 1790.8538533533533u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1794.7630135135132u,0 1794.7640135135134u,1.5 1795.7405535535534u,1.5 1795.7415535535536u,0 1802.5833338338336u,0 1802.5843338338339u,1.5 1803.5608738738738u,1.5 1803.561873873874u,0 1804.5384139139137u,0 1804.539413913914u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1823.1116746746745u,0 1823.1126746746747u,1.5 1824.0892147147147u,1.5 1824.0902147147149u,0 1826.0442947947947u,0 1826.045294794795u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1839.7298553553553u,1.5 1839.7308553553555u,0 1851.4603358358356u,0 1851.4613358358358u,1.5 1855.370495995996u,1.5 1855.3714959959962u,0 1856.3480360360359u,0 1856.349036036036u,1.5 1863.1908163163164u,1.5 1863.1918163163166u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1866.1234364364361u,1.5 1866.1244364364363u,0 1876.8763768768767u,0 1876.877376876877u,1.5 1877.853916916917u,1.5 1877.854916916917u,0 1878.8314569569568u,0 1878.832456956957u,1.5 1889.5843973973974u,1.5 1889.5853973973976u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1896.4271776776775u,1.5 1896.4281776776777u,0 1897.4047177177176u,0 1897.4057177177178u,1.5 1898.3822577577575u,1.5 1898.3832577577577u,0 1899.3597977977977u,0 1899.3607977977979u,1.5 1900.3373378378376u,1.5 1900.3383378378378u,0 1911.0902782782782u,0 1911.0912782782784u,1.5 1915.0004384384383u,1.5 1915.0014384384385u,0 1916.9555185185184u,0 1916.9565185185186u,1.5 1929.6635390390388u,1.5 1929.664539039039u,0 1930.641079079079u,0 1930.6420790790792u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1940.4164794794794u,0 1940.4174794794797u,1.5 1941.3940195195194u,1.5 1941.3950195195196u,0 1943.3490995995994u,0 1943.3500995995996u,1.5 1944.3266396396396u,1.5 1944.3276396396398u,0 1958.9897402402403u,0 1958.9907402402405u,1.5 1959.9672802802804u,1.5 1959.9682802802806u,0 1960.94482032032u,0 1960.9458203203203u,1.5 1961.9223603603602u,1.5 1961.9233603603604u,0 1964.8549804804804u,0 1964.8559804804806u,1.5 1965.8325205205203u,1.5 1965.8335205205206u,0 1967.7876006006004u,0 1967.7886006006006u,1.5 1968.7651406406405u,1.5 1968.7661406406407u,0 1970.7202207207204u,0 1970.7212207207206u,1.5 1971.6977607607605u,1.5 1971.6987607607607u,0 1974.630380880881u,0 1974.6313808808811u,1.5 1976.5854609609607u,1.5 1976.586460960961u,0 1977.5630010010009u,0 1977.564001001001u,1.5 1980.4956211211208u,1.5 1980.496621121121u,0 1981.473161161161u,0 1981.4741611611612u,1.5 1983.4282412412413u,1.5 1983.4292412412415u,0 1984.4057812812814u,0 1984.4067812812816u,1.5 1987.3384014014014u,1.5 1987.3394014014016u,0 1988.3159414414415u,0 1988.3169414414417u,1.5 1989.2934814814816u,1.5 1989.2944814814819u,0 1990.2710215215213u,0 1990.2720215215215u,1.5 1995.1587217217213u,1.5 1995.1597217217216u,0 1996.1362617617615u,0 1996.1372617617617u,1.5 1998.0913418418418u,1.5 1998.092341841842u,0 1999.068881881882u,0 1999.069881881882u,1.5 2007.8667422422423u,1.5 2007.8677422422425u,0 2008.8442822822824u,0 2008.8452822822826u,1.5 2014.7095225225223u,1.5 2014.7105225225225u,0 2015.6870625625625u,0 2015.6880625625627u,1.5 2021.5523028028026u,1.5 2021.5533028028028u,0 2022.5298428428428u,0 2022.530842842843u,1.5 2023.507382882883u,1.5 2023.508382882883u,0 2024.4849229229226u,0 2024.4859229229228u,1.5 2025.4624629629627u,1.5 2025.463462962963u,0 2026.4400030030029u,0 2026.441003003003u,1.5 2027.417543043043u,1.5 2027.4185430430432u,0 2028.3950830830831u,0 2028.3960830830833u,1.5 2029.3726231231228u,1.5 2029.373623123123u,0 2032.3052432432432u,0 2032.3062432432434u,1.5 2033.2827832832834u,1.5 2033.2837832832836u,0 2036.2154034034033u,0 2036.2164034034035u,1.5 2037.1929434434435u,1.5 2037.1939434434437u,0 2041.1031036036034u,0 2041.1041036036036u,1.5 2042.0806436436435u,1.5 2042.0816436436437u,0 2059.676364364364u,0 2059.677364364364u,1.5 2060.6539044044043u,1.5 2060.6549044044045u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2067.4966846846846u,0 2067.497684684685u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2070.429304804805u,0 2070.430304804805u,1.5 2086.0699454454452u,1.5 2086.0709454454454u,0 2091.9351856856856u,0 2091.936185685686u,1.5 2092.9127257257255u,1.5 2092.9137257257257u,0 2103.665666166166u,0 2103.666666166166u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2105.620746246246u,0 2105.6217462462464u,1.5 2120.2838468468467u,1.5 2120.284846846847u,0 2121.261386886887u,0 2121.2623868868873u,1.5 2123.216466966967u,1.5 2123.217466966967u,0 2134.946947447447u,0 2134.9479474474474u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2137.8795675675674u,0 2137.8805675675676u,1.5 2138.8571076076073u,1.5 2138.8581076076075u,0 2139.8346476476477u,0 2139.835647647648u,1.5 2149.610048048048u,1.5 2149.6110480480484u,0 2162.3180685685684u,0 2162.3190685685686u,1.5 2163.2956086086083u,1.5 2163.2966086086085u,0 2164.2731486486487u,0 2164.274148648649u,1.5 2174.048549049049u,1.5 2174.0495490490493u,0 2184.8014894894895u,0 2184.8024894894897u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2187.7341096096093u,0 2187.7351096096095u,1.5 2196.53196996997u,1.5 2196.53296996997u,0 2197.5095100100098u,0 2197.51051001001u,1.5 2198.48705005005u,1.5 2198.4880500500503u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2219.992930930931u,1.5 2219.993930930931u,0 2220.970470970971u,0 2220.971470970971u,1.5 2221.9480110110107u,1.5 2221.949011011011u,0 2227.813251251251u,0 2227.8142512512513u,1.5 2228.790791291291u,1.5 2228.7917912912912u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2230.745871371371u,1.5 2230.746871371371u,0 2231.7234114114112u,0 2231.7244114114114u,1.5 2238.5661916916915u,1.5 2238.5671916916917u,0 2239.543731731732u,0 2239.544731731732u,1.5 2240.5212717717714u,1.5 2240.5222717717716u,0 2241.4988118118117u,0 2241.499811811812u,1.5 2242.4763518518516u,1.5 2242.477351851852u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2254.2068323323324u,0 2254.2078323323326u,1.5 2260.0720725725723u,1.5 2260.0730725725725u,0 2268.869932932933u,0 2268.870932932933u,1.5 2269.847472972973u,1.5 2269.848472972973u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2280.600413413413u,1.5 2280.6014134134134u,0 2281.577953453453u,0 2281.5789534534533u,1.5 2282.5554934934935u,1.5 2282.5564934934937u,0 2290.3758138138137u,0 2290.376813813814u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2293.308433933934u,0 2293.309433933934u,1.5 2304.0613743743743u,1.5 2304.0623743743745u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2314.8143148148147u,1.5 2314.815314814815u,0 2316.769394894895u,0 2316.770394894895u,1.5 2317.746934934935u,1.5 2317.747934934935u,0 2318.724474974975u,0 2318.725474974975u,1.5 2324.589715215215u,1.5 2324.5907152152154u,0 2325.567255255255u,0 2325.5682552552553u,1.5 2327.5223353353354u,1.5 2327.5233353353356u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2340.2303558558556u,1.5 2340.231355855856u,0 2341.207895895896u,0 2341.208895895896u,1.5 2349.028216216216u,1.5 2349.0292162162164u,0 2350.005756256256u,0 2350.0067562562563u,1.5 2350.9832962962964u,1.5 2350.9842962962966u,0 2359.7811566566565u,0 2359.7821566566568u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2365.646396896897u,0 2365.647396896897u,1.5 2367.6014769769768u,1.5 2367.602476976977u,0 2368.5790170170167u,0 2368.580017017017u,1.5 2376.3993373373373u,1.5 2376.4003373373375u,0 2377.3768773773777u,0 2377.377877377378u,1.5 2380.3094974974974u,1.5 2380.3104974974976u,0 2393.995058058058u,0 2393.996058058058u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2397.905218218218u,0 2397.9062182182183u,1.5 2410.613238738739u,1.5 2410.614238738739u,0 2411.5907787787787u,0 2411.591778778779u,1.5 2412.5683188188186u,1.5 2412.569318818819u,0 2415.500938938939u,0 2415.501938938939u,1.5 2416.478478978979u,1.5 2416.4794789789794u,0 2432.119119619619u,0 2432.1201196196193u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2435.05173973974u,1.5 2435.05273973974u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.9843598598595u,1.5 2437.9853598598597u,0 2438.9618998999u,0 2438.9628998999u,1.5 2459.490240740741u,1.5 2459.491240740741u,0 2460.4677807807807u,0 2460.468780780781u,1.5 2461.4453208208206u,1.5 2461.446320820821u,0 2462.4228608608605u,0 2462.4238608608607u,1.5 2464.377940940941u,1.5 2464.378940940941u,0 2465.355480980981u,0 2465.3564809809814u,1.5 2466.3330210210206u,1.5 2466.334021021021u,0 2467.310561061061u,0 2467.311561061061u,1.5 2468.288101101101u,1.5 2468.289101101101u,0 2472.198261261261u,0 2472.199261261261u,1.5 2474.1533413413413u,1.5 2474.1543413413415u,0 2476.108421421421u,0 2476.1094214214213u,1.5 2478.0635015015014u,1.5 2478.0645015015016u,0 2482.9512017017014u,0 2482.9522017017016u,1.5 2483.9287417417418u,1.5 2483.929741741742u,0 2484.9062817817817u,0 2484.907281781782u,1.5 2485.8838218218216u,1.5 2485.884821821822u,0 2501.5244624624625u,0 2501.5254624624627u,1.5 2502.5020025025024u,1.5 2502.5030025025026u,0 2503.4795425425427u,0 2503.480542542543u,1.5 2504.4570825825826u,1.5 2504.458082582583u,0 2512.277402902903u,0 2512.278402902903u,1.5 2513.2549429429428u,1.5 2513.255942942943u,0 2517.165103103103u,0 2517.166103103103u,1.5 2518.1426431431432u,1.5 2518.1436431431434u,0 2519.120183183183u,0 2519.1211831831833u,1.5 2520.097723223223u,1.5 2520.0987232232233u,0 2522.0528033033033u,0 2522.0538033033035u,1.5 2523.0303433433432u,1.5 2523.0313433433435u,0 2524.985423423423u,0 2524.9864234234233u,1.5 2525.9629634634634u,1.5 2525.9639634634636u,0 2527.9180435435437u,0 2527.919043543544u,1.5 2528.8955835835836u,1.5 2528.896583583584u,0 2529.8731236236235u,0 2529.8741236236237u,1.5 2531.8282037037034u,1.5 2531.8292037037036u,0 2532.8057437437437u,0 2532.806743743744u,1.5 2533.7832837837836u,1.5 2533.784283783784u,0 2534.7608238238236u,0 2534.7618238238238u,1.5 2544.536224224224u,1.5 2544.5372242242242u,0 2545.513764264264u,0 2545.514764264264u,1.5 2554.3116246246245u,1.5 2554.3126246246247u,0 2555.2891646646644u,0 2555.2901646646646u,1.5 2558.2217847847846u,1.5 2558.222784784785u,0 2559.1993248248245u,0 2559.2003248248247u,1.5 2560.1768648648645u,1.5 2560.1778648648647u,0 2562.1319449449447u,0 2562.132944944945u,1.5 2565.064565065065u,1.5 2565.065565065065u,0 2566.042105105105u,0 2566.043105105105u,1.5 2567.019645145145u,1.5 2567.0206451451454u,0 2567.997185185185u,0 2567.9981851851853u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2586.5704459459457u,0 2586.571445945946u,1.5 2587.547985985986u,1.5 2587.5489859859863u,0 2588.5255260260255u,0 2588.5265260260257u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2608.0763268268265u,1.5 2608.0773268268267u,0 2619.8068073073073u,0 2619.8078073073075u,1.5 2620.784347347347u,1.5 2620.7853473473474u,0 2622.739427427427u,0 2622.740427427427u,1.5 2634.469907907908u,1.5 2634.470907907908u,0 2635.4474479479477u,0 2635.448447947948u,1.5 2637.402528028028u,1.5 2637.403528028028u,0 2650.1105485485486u,0 2650.111548548549u,1.5 2652.065628628629u,1.5 2652.066628628629u,0 2653.0431686686684u,0 2653.0441686686686u,1.5 2657.9308688688684u,1.5 2657.9318688688686u,0 2658.9084089089088u,0 2658.909408908909u,1.5 2659.8859489489487u,1.5 2659.886948948949u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2665.751189189189u,0 2665.7521891891893u,1.5 2666.7287292292294u,1.5 2666.7297292292296u,0 2672.5939694694694u,0 2672.5949694694696u,1.5 2673.5715095095093u,1.5 2673.5725095095095u,0 2674.5490495495496u,0 2674.55004954955u,1.5 2685.30198998999u,1.5 2685.3029899899902u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2689.21215015015u,0 2689.2131501501503u,1.5 2690.18969019019u,1.5 2690.1906901901903u,0 2694.09985035035u,0 2694.1008503503504u,1.5 2695.0773903903905u,1.5 2695.0783903903907u,0 2696.0549304304304u,0 2696.0559304304306u,1.5 2698.0100105105103u,1.5 2698.0110105105105u,0 2698.9875505505506u,0 2698.988550550551u,1.5 2699.9650905905905u,1.5 2699.9660905905907u,0 2700.942630630631u,0 2700.943630630631u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2710.718031031031u,0 2710.719031031031u,1.5 2711.695571071071u,1.5 2711.696571071071u,0 2718.538351351351u,0 2718.5393513513513u,1.5 2719.5158913913915u,1.5 2719.5168913913917u,0 2720.4934314314314u,0 2720.4944314314316u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2730.268831831832u,1.5 2730.269831831832u,0 2737.1116121121117u,0 2737.112612112112u,1.5 2738.089152152152u,1.5 2738.0901521521523u,0 2739.066692192192u,0 2739.067692192192u,1.5 2740.0442322322324u,1.5 2740.0452322322326u,0 2741.021772272272u,0 2741.022772272272u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2750.7971726726723u,1.5 2750.7981726726725u,0 2751.7747127127127u,0 2751.775712712713u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 2756.6624129129127u,0 2756.663412912913u,1.5 2757.6399529529526u,1.5 2757.640952952953u,0 2760.572573073073u,0 2760.573573073073u,1.5 2761.5501131131127u,1.5 2761.551113113113u,0 2762.527653153153u,0 2762.5286531531533u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2773.2805935935935u,1.5 2773.2815935935937u,0 2782.0784539539536u,0 2782.079453953954u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2801.6292547547546u,0 2801.630254754755u,1.5 2803.584334834835u,1.5 2803.585334834835u,0 2804.561874874875u,0 2804.562874874875u,1.5 2805.5394149149147u,1.5 2805.540414914915u,0 2806.5169549549546u,0 2806.517954954955u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2822.1575955955955u,0 2822.1585955955957u,1.5 2823.135135635636u,1.5 2823.136135635636u,0 2824.1126756756753u,0 2824.1136756756755u,1.5 2825.0902157157157u,1.5 2825.091215715716u,0 2826.0677557557556u,0 2826.068755755756u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2839.753316316316u,0 2839.7543163163164u,1.5 2840.730856356356u,1.5 2840.7318563563563u,0 2848.5511766766763u,0 2848.5521766766765u,1.5 2850.5062567567566u,1.5 2850.5072567567568u,0 2852.461336836837u,0 2852.462336836837u,1.5 2860.281657157157u,1.5 2860.2826571571572u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2865.169357357357u,0 2865.1703573573573u,1.5 2866.1468973973974u,1.5 2866.1478973973976u,0 2875.922297797798u,0 2875.923297797798u,1.5 2876.899837837838u,1.5 2876.900837837838u,0 2877.877377877878u,0 2877.8783778778784u,1.5 2878.8549179179176u,1.5 2878.855917917918u,0 2879.832457957958u,0 2879.833457957958u,1.5 2880.809997997998u,1.5 2880.810997997998u,0 2881.787538038038u,0 2881.788538038038u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2909.158659159159u,0 2909.159659159159u,1.5 2910.136199199199u,1.5 2910.137199199199u,0 2912.091279279279u,0 2912.0922792792794u,1.5 2913.068819319319u,1.5 2913.0698193193193u,0 2914.046359359359u,0 2914.0473593593592u,1.5 2930.66454004004u,1.5 2930.66554004004u,0 2931.64208008008u,0 2931.6430800800804u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2938.48486036036u,0 2938.48586036036u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2941.4174804804807u,1.5 2941.418480480481u,0 2942.39502052052u,0 2942.3960205205203u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 2958.035661161161u,0 2958.036661161161u,1.5 2959.013201201201u,1.5 2959.014201201201u,0 2962.923361361361u,0 2962.924361361361u,1.5 2963.9009014014014u,1.5 2963.9019014014016u,0 2965.8559814814816u,0 2965.856981481482u,1.5 2966.833521521521u,1.5 2966.8345215215213u,0 2968.7886016016014u,0 2968.7896016016016u,1.5 2969.7661416416418u,1.5 2969.767141641642u,0 2970.7436816816817u,0 2970.744681681682u,1.5 2971.7212217217216u,1.5 2971.722221721722u,0 2972.6987617617615u,0 2972.6997617617617u,1.5 2973.676301801802u,1.5 2973.677301801802u,0 2974.6538418418418u,0 2974.654841841842u,1.5 2979.541542042042u,1.5 2979.542542042042u,0 2980.519082082082u,0 2980.5200820820824u,1.5 2982.474162162162u,1.5 2982.475162162162u,0 2983.451702202202u,0 2983.452702202202u,1.5 2992.2495625625625u,1.5 2992.2505625625627u,0 2993.2271026026024u,0 2993.2281026026026u,1.5 3006.912663163163u,1.5 3006.913663163163u,0 3007.890203203203u,0 3007.891203203203u,1.5 3008.8677432432432u,1.5 3008.8687432432434u,0 3009.845283283283u,0 3009.8462832832834u,1.5 3010.822823323323u,1.5 3010.8238233233233u,0 3011.800363363363u,0 3011.801363363363u,1.5 3013.7554434434433u,1.5 3013.7564434434435u,0 3014.7329834834836u,0 3014.733983483484u,1.5 3016.6880635635634u,1.5 3016.6890635635636u,0 3017.6656036036034u,0 3017.6666036036036u,1.5 3018.6431436436437u,1.5 3018.644143643644u,0 3019.6206836836836u,0 3019.621683683684u,1.5 3022.553303803804u,1.5 3022.554303803804u,0 3024.508383883884u,0 3024.5093838838843u,1.5 3025.4859239239236u,1.5 3025.4869239239238u,0 3027.441004004004u,0 3027.442004004004u,1.5 3028.418544044044u,1.5 3028.4195440440444u,0 3029.396084084084u,0 3029.3970840840843u,1.5 3030.373624124124u,1.5 3030.3746241241242u,0 3032.328704204204u,0 3032.329704204204u,1.5 3033.306244244244u,1.5 3033.3072442442444u,0 3034.283784284284u,0 3034.2847842842843u,1.5 3035.261324324324u,1.5 3035.2623243243243u,0 3038.1939444444442u,0 3038.1949444444444u,1.5 3039.1714844844846u,1.5 3039.172484484485u,0 3042.1041046046043u,0 3042.1051046046045u,1.5 3043.0816446446447u,1.5 3043.082644644645u,0 3062.6324454454452u,0 3062.6334454454454u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3066.5426056056053u,1.5 3066.5436056056055u,0 3067.5201456456457u,0 3067.521145645646u,1.5 3084.138326326326u,1.5 3084.139326326326u,0 3085.115866366366u,0 3085.116866366366u,1.5 3088.0484864864866u,1.5 3088.049486486487u,0 3090.0035665665664u,0 3090.0045665665666u,1.5 3090.9811066066063u,1.5 3090.9821066066065u,0 3103.689127127127u,0 3103.690127127127u,1.5 3104.666667167167u,1.5 3104.667667167167u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3118.3522277277275u,1.5 3118.3532277277277u,0 3120.307307807808u,0 3120.308307807808u,1.5 3122.262387887888u,1.5 3122.2633878878883u,0 3125.195008008008u,0 3125.196008008008u,1.5 3126.172548048048u,1.5 3126.1735480480484u,0 3135.947948448448u,0 3135.9489484484484u,1.5 3147.678428928929u,1.5 3147.679428928929u,0 3148.655968968969u,0 3148.656968968969u,1.5 3151.588589089089u,1.5 3151.5895890890893u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3175.04955005005u,1.5 3175.0505500500503u,0 3177.0046301301304u,0 3177.0056301301306u,1.5 3177.98217017017u,1.5 3177.98317017017u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3196.555430930931u,1.5 3196.556430930931u,0 3197.532970970971u,0 3197.533970970971u,1.5 3198.5105110110107u,1.5 3198.511511011011u,0 3207.308371371371u,0 3207.309371371371u,1.5 3216.106231731732u,1.5 3216.107231731732u,0 3217.0837717717714u,0 3217.0847717717716u,1.5 3218.0613118118117u,1.5 3218.062311811812u,0 3219.0388518518516u,0 3219.039851851852u,1.5 3220.016391891892u,1.5 3220.017391891892u,0 3227.836712212212u,0 3227.8377122122124u,1.5 3228.814252252252u,1.5 3228.8152522522523u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3232.724412412412u,1.5 3232.7254124124124u,0 3233.701952452452u,0 3233.7029524524523u,1.5 3237.6121126126122u,1.5 3237.6131126126124u,0 3238.5896526526526u,0 3238.590652652653u,1.5 3239.5671926926925u,1.5 3239.5681926926927u,0 3240.544732732733u,0 3240.545732732733u,1.5 3241.5222727727723u,1.5 3241.5232727727725u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3259.1179934934935u,1.5 3259.1189934934937u,0 3260.0955335335334u,0 3260.0965335335336u,1.5 3262.050613613613u,1.5 3262.0516136136134u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3273.781094094094u,0 3273.782094094094u,1.5 3278.6687942942945u,1.5 3278.6697942942947u,0 3279.6463343343344u,0 3279.6473343343346u,1.5 3280.6238743743743u,1.5 3280.6248743743745u,0 3281.601414414414u,0 3281.6024144144144u,1.5 3283.5564944944945u,1.5 3283.5574944944947u,0 3290.3992747747743u,0 3290.4002747747745u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3294.309434934935u,0 3294.310434934935u,1.5 3302.129755255255u,1.5 3302.1307552552553u,0 3303.1072952952954u,0 3303.1082952952956u,1.5 3304.0848353353354u,1.5 3304.0858353353356u,0 3309.9500755755753u,0 3309.9510755755755u,1.5 3310.927615615615u,1.5 3310.9286156156154u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3325.590716216216u,1.5 3325.5917162162164u,0 3335.366116616616u,0 3335.3671166166164u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3349.0516771771768u,1.5 3349.052677177177u,0 3350.029217217217u,0 3350.0302172172173u,1.5 3351.006757257257u,1.5 3351.0077572572573u,0 3351.9842972972974u,0 3351.9852972972976u,1.5 3352.9618373373373u,1.5 3352.9628373373375u,0 3353.9393773773772u,0 3353.9403773773774u,1.5 3354.916917417417u,1.5 3354.9179174174174u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3365.6698578578576u,1.5 3365.6708578578578u,0 3366.647397897898u,0 3366.648397897898u,1.5 3378.3778783783787u,1.5 3378.378878378379u,0 3383.2655785785787u,0 3383.266578578579u,1.5 3384.243118618618u,1.5 3384.2441186186184u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3390.1083588588585u,1.5 3390.1093588588587u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3396.9511391391393u,0 3396.9521391391395u,1.5 3409.6591596596595u,1.5 3409.6601596596597u,0 3410.6366996996994u,0 3410.6376996996996u,1.5 3413.5693198198196u,1.5 3413.57031981982u,0 3415.5243998999u,0 3415.5253998999u,1.5 3417.47947997998u,1.5 3417.4804799799804u,0 3418.4570200200196u,0 3418.45802002002u,1.5 3419.43456006006u,1.5 3419.43556006006u,0 3431.1650405405403u,0 3431.1660405405405u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3434.0976606606605u,0 3434.0986606606607u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3436.052740740741u,0 3436.053740740741u,1.5 3455.6035415415413u,1.5 3455.6045415415415u,0 3456.5810815815817u,0 3456.582081581582u,1.5 3458.5361616616615u,1.5 3458.5371616616617u,0 3459.5137017017014u,0 3459.5147017017016u,1.5 3463.4238618618615u,1.5 3463.4248618618617u,0 3464.401401901902u,0 3464.402401901902u,1.5 3466.356481981982u,1.5 3466.3574819819823u,0 3468.311562062062u,0 3468.312562062062u,1.5 3469.289102102102u,1.5 3469.290102102102u,0 3471.244182182182u,0 3471.2451821821824u,1.5 3472.221722222222u,1.5 3472.2227222222223u,0 3475.1543423423423u,0 3475.1553423423425u,1.5 3476.1318823823826u,1.5 3476.132882382383u,0 3478.0869624624625u,0 3478.0879624624627u,1.5 3479.0645025025024u,1.5 3479.0655025025026u,0 3484.9297427427427u,0 3484.930742742743u,1.5 3485.9072827827827u,1.5 3485.908282782783u,0 3486.8848228228226u,0 3486.885822822823u,1.5 3487.8623628628625u,1.5 3487.8633628628627u,0 3488.839902902903u,0 3488.840902902903u,1.5 3489.8174429429428u,1.5 3489.818442942943u,0 3497.637763263263u,0 3497.638763263263u,1.5 3498.6153033033033u,1.5 3498.6163033033035u,0 3500.5703833833836u,0 3500.571383383384u,1.5 3501.547923423423u,1.5 3501.5489234234233u,0 3511.3233238238236u,0 3511.3243238238238u,1.5 3512.3008638638635u,1.5 3512.3018638638637u,0 3514.2559439439437u,0 3514.256943943944u,1.5 3515.233483983984u,1.5 3515.2344839839843u,0 3521.098724224224u,0 3521.0997242242242u,1.5 3522.076264264264u,1.5 3522.077264264264u,0 3524.0313443443442u,0 3524.0323443443444u,1.5 3525.986424424424u,1.5 3525.9874244244243u,0 3527.9415045045043u,0 3527.9425045045045u,1.5 3528.9190445445447u,1.5 3528.920044544545u,0 3529.8965845845846u,0 3529.897584584585u,1.5 3530.8741246246245u,1.5 3530.8751246246247u,0 3532.8292047047044u,0 3532.8302047047046u,1.5 3538.6944449449447u,1.5 3538.695444944945u,0 3539.671984984985u,0 3539.6729849849853u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.020646146146u,0 3568.0216461461464u,1.5 3568.998186186186u,1.5 3568.9991861861863u,0 3577.7960465465467u,0 3577.797046546547u,1.5 3578.7735865865866u,1.5 3578.774586586587u,0 3586.593906906907u,0 3586.594906906907u,1.5 3587.5714469469467u,1.5 3587.572446946947u,0 3588.548986986987u,0 3588.5499869869873u,1.5 3591.481607107107u,1.5 3591.482607107107u,0 3592.459147147147u,0 3592.4601471471474u,1.5 3603.2120875875876u,1.5 3603.213087587588u,0 3605.1671676676674u,0 3605.1681676676676u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3607.1222477477477u,0 3607.123247747748u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3621.785348348348u,0 3621.7863483483484u,1.5 3623.740428428428u,1.5 3623.741428428428u,0 3624.7179684684684u,0 3624.7189684684686u,1.5 3635.4709089089088u,1.5 3635.471908908909u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3637.425988988989u,1.5 3637.4269889889893u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3646.223849349349u,0 3646.2248493493494u,1.5 3647.2013893893895u,1.5 3647.2023893893897u,0 3651.1115495495496u,0 3651.11254954955u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3673.5949704704703u,0 3673.5959704704705u,1.5 3674.5725105105103u,1.5 3674.5735105105105u,0 3675.5500505505506u,0 3675.551050550551u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3688.258071071071u,1.5 3688.259071071071u,0 3697.0559314314314u,0 3697.0569314314316u,1.5 3699.9885515515516u,1.5 3699.989551551552u,0 3700.9660915915915u,0 3700.9670915915917u,1.5 3706.831331831832u,1.5 3706.832331831832u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3717.584272272272u,0 3717.585272272272u,1.5 3719.539352352352u,1.5 3719.5403523523523u,0 3720.5168923923925u,0 3720.5178923923927u,1.5 3721.4944324324324u,1.5 3721.4954324324326u,0 3722.4719724724723u,0 3722.4729724724725u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3732.2473728728723u,0 3732.2483728728726u,1.5 3733.2249129129127u,1.5 3733.225912912913u,0 3739.090153153153u,0 3739.0911531531533u,1.5 3740.067693193193u,1.5 3740.068693193193u,0 3741.0452332332334u,0 3741.0462332332336u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3757.6634139139137u,0 3757.664413913914u,1.5 3758.6409539539536u,1.5 3758.641953953954u,0 3759.618493993994u,0 3759.619493993994u,1.5 3760.596034034034u,1.5 3760.597034034034u,0 3761.573574074074u,0 3761.574574074074u,1.5 3772.326514514514u,1.5 3772.3275145145144u,0 3780.146834834835u,0 3780.147834834835u,1.5 3781.124374874875u,1.5 3781.125374874875u,0 3783.0794549549546u,0 3783.080454954955u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3802.6302557557556u,0 3802.631255755756u,1.5 3803.607795795796u,1.5 3803.608795795796u,0 3804.585335835836u,0 3804.586335835836u,1.5 3806.5404159159157u,1.5 3806.541415915916u,0 3807.5179559559556u,0 3807.518955955956u,1.5 3812.405656156156u,1.5 3812.4066561561563u,0 3813.383196196196u,0 3813.384196196196u,1.5 3814.3607362362363u,1.5 3814.3617362362365u,0 3815.338276276276u,0 3815.339276276276u,1.5 3816.315816316316u,1.5 3816.3168163163164u,0 3817.293356356356u,0 3817.2943563563563u,1.5 3818.2708963963964u,1.5 3818.2718963963966u,0 3825.1136766766763u,0 3825.1146766766765u,1.5 3826.0912167167166u,1.5 3826.092216716717u,0 3827.0687567567566u,0 3827.0697567567568u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3836.844157157157u,0 3836.8451571571572u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 3847.5970975975974u,0 3847.5980975975976u,1.5 3848.574637637638u,1.5 3848.575637637638u,0 3850.5297177177176u,0 3850.530717717718u,1.5 3851.5072577577575u,1.5 3851.5082577577577u,0 3852.484797797798u,0 3852.485797797798u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3876.923298798799u,0 3876.924298798799u,1.5 3877.900838838839u,1.5 3877.901838838839u,0 3879.8559189189186u,0 3879.856918918919u,1.5 3887.6762392392393u,1.5 3887.6772392392395u,0 3888.653779279279u,0 3888.6547792792794u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3895.4965595595595u,1.5 3895.4975595595597u,0 3913.09228028028u,0 3913.0932802802804u,1.5 3914.06982032032u,1.5 3914.0708203203203u,0 3915.0473603603605u,0 3915.0483603603607u,1.5 3917.00244044044u,1.5 3917.00344044044u,0 3917.9799804804807u,0 3917.980980480481u,1.5 3933.6206211211206u,1.5 3933.621621121121u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3938.508321321321u,0 3938.5093213213213u,1.5 3939.4858613613615u,1.5 3939.4868613613617u,0 3960.991742242242u,0 3960.992742242242u,1.5 3961.969282282282u,1.5 3961.9702822822824u,0 3962.946822322322u,0 3962.9478223223223u,1.5 3963.9243623623624u,1.5 3963.9253623623626u,0 3965.879442442442u,0 3965.880442442442u,1.5 3966.8569824824826u,1.5 3966.857982482483u,0 3967.834522522522u,0 3967.8355225225223u,1.5 3969.7896026026024u,1.5 3969.7906026026026u,0 3972.7222227227226u,0 3972.7232227227228u,1.5 3973.699762762763u,1.5 3973.700762762763u,0 3974.677302802803u,0 3974.678302802803u,1.5 3975.6548428428423u,1.5 3975.6558428428425u,0 3977.6099229229226u,0 3977.610922922923u,1.5 3980.5425430430428u,1.5 3980.543543043043u,0 3981.520083083083u,0 3981.5210830830833u,1.5 3982.4976231231226u,1.5 3982.498623123123u,0 3983.4751631631634u,0 3983.4761631631636u,1.5 3989.3404034034033u,1.5 3989.3414034034035u,0 3990.317943443443u,0 3990.318943443443u,1.5 3998.138263763764u,1.5 3998.139263763764u,0 3999.115803803804u,0 3999.116803803804u,1.5 4013.7789044044043u,1.5 4013.7799044044045u,0 4014.756444444444u,0 4014.757444444444u,1.5 4016.711524524524u,1.5 4016.7125245245243u,0 4017.689064564565u,0 4017.690064564565u,1.5 4020.6216846846846u,1.5 4020.622684684685u,0 4021.5992247247245u,0 4021.6002247247247u,1.5 4024.5318448448443u,1.5 4024.5328448448445u,0 4026.4869249249246u,0 4026.4879249249248u,1.5 4027.4644649649654u,1.5 4027.4654649649656u,0 4028.442005005005u,0 4028.443005005005u,1.5 4029.4195450450447u,1.5 4029.420545045045u,0 4030.397085085085u,0 4030.3980850850853u,1.5 4031.374625125125u,1.5 4031.375625125125u,0 4033.329705205205u,0 4033.330705205205u,1.5 4035.284785285285u,1.5 4035.2857852852853u,0 4037.2398653653654u,0 4037.2408653653656u,1.5 4038.2174054054053u,1.5 4038.2184054054055u,0 4039.194945445445u,0 4039.195945445445u,1.5 4040.1724854854856u,1.5 4040.173485485486u,0 4043.1051056056053u,0 4043.1061056056055u,1.5 4044.0826456456452u,1.5 4044.0836456456454u,0 4057.768206206206u,0 4057.769206206206u,1.5 4058.7457462462457u,1.5 4058.746746246246u,0 4061.6783663663664u,0 4061.6793663663666u,1.5 4062.6559064064063u,1.5 4062.6569064064065u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4065.588526526526u,1.5 4065.5895265265262u,0 4066.566066566567u,0 4066.567066566567u,1.5 4067.5436066066063u,1.5 4067.5446066066065u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4080.251627127127u,1.5 4080.252627127127u,0 4081.2291671671674u,0 4081.2301671671676u,1.5 4084.161787287287u,1.5 4084.1627872872873u,0 4085.139327327327u,0 4085.140327327327u,1.5 4086.1168673673674u,1.5 4086.1178673673676u,0 4087.0944074074073u,0 4087.0954074074075u,1.5 4089.0494874874876u,1.5 4089.0504874874878u,0 4093.9371876876876u,0 4093.938187687688u,1.5 4094.9147277277275u,1.5 4094.9157277277277u,0 4101.757508008008u,0 4101.758508008008u,1.5 4102.735048048047u,1.5 4102.736048048047u,0 4104.690128128128u,0 4104.691128128128u,1.5 4105.667668168168u,1.5 4105.668668168169u,0 4106.645208208208u,0 4106.646208208208u,1.5 4119.353228728728u,1.5 4119.354228728728u,0 4120.330768768769u,0 4120.3317687687695u,1.5 4122.285848848848u,1.5 4122.286848848848u,0 4124.240928928929u,0 4124.241928928929u,1.5 4125.218468968969u,1.5 4125.2194689689695u,0 4134.993869369369u,0 4134.99486936937u,1.5 4137.9264894894895u,1.5 4137.92748948949u,0 4138.904029529529u,0 4138.905029529529u,1.5 4146.724349849849u,1.5 4146.725349849849u,0 4147.70188988989u,0 4147.70288988989u,1.5 4148.67942992993u,1.5 4148.68042992993u,0 4149.65696996997u,0 4149.6579699699705u,1.5 4150.63451001001u,1.5 4150.63551001001u,0 4161.38745045045u,0 4161.38845045045u,1.5 4172.140390890891u,1.5 4172.141390890891u,0 4173.117930930931u,0 4173.118930930931u,1.5 4174.095470970971u,1.5 4174.0964709709715u,0 4183.870871371371u,0 4183.8718713713715u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4193.646271771772u,1.5 4193.6472717717725u,0 4194.623811811812u,0 4194.624811811812u,1.5 4197.556431931932u,1.5 4197.557431931932u,0 4198.533971971972u,0 4198.5349719719725u,1.5 4199.511512012012u,1.5 4199.512512012012u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4209.286912412412u,0 4209.287912412412u,1.5 4219.062312812813u,1.5 4219.063312812813u,0 4225.9050930930935u,0 4225.906093093094u,1.5 4226.882633133133u,1.5 4226.883633133133u,0 4229.815253253253u,0 4229.816253253253u,1.5 4236.658033533533u,1.5 4236.659033533533u,0 4237.635573573573u,0 4237.6365735735735u,1.5 4238.613113613614u,1.5 4238.614113613614u,0 4239.590653653653u,0 4239.591653653653u,1.5 4240.5681936936935u,1.5 4240.569193693694u,0 4251.321134134134u,0 4251.322134134134u,1.5 4260.1189944944945u,1.5 4260.119994494495u,0 4261.096534534534u,0 4261.097534534534u,1.5 4262.074074574574u,1.5 4262.0750745745745u,0 4268.916854854855u,0 4268.917854854855u,1.5 4270.871934934935u,1.5 4270.872934934935u,0 4272.827015015015u,0 4272.828015015015u,1.5 4282.602415415415u,1.5 4282.603415415415u,0 4289.4451956956955u,0 4289.446195695696u,1.5 4290.422735735735u,1.5 4290.423735735735u,0 4292.377815815816u,0 4292.378815815816u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4294.3328958958955u,0 4294.333895895896u,1.5 4303.130756256257u,1.5 4303.131756256257u,0 4313.8836966966965u,0 4313.884696696697u,1.5 4322.681557057057u,1.5 4322.682557057057u,0 4323.659097097097u,0 4323.660097097098u,1.5 4326.591717217217u,1.5 4326.592717217217u,0 4327.569257257258u,0 4327.570257257258u,1.5 4328.546797297297u,1.5 4328.547797297298u,0 4336.367117617618u,0 4336.368117617618u,1.5 4337.344657657658u,1.5 4337.345657657658u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4342.232357857858u,0 4342.233357857858u,1.5 4347.120058058058u,1.5 4347.121058058058u,0 4348.097598098098u,0 4348.098598098099u,1.5 4351.030218218218u,1.5 4351.031218218218u,0 4361.783158658659u,0 4361.784158658659u,1.5 4362.760698698698u,1.5 4362.761698698699u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4368.625938938939u,1.5 4368.626938938939u,0 4369.603478978979u,0 4369.604478978979u,1.5 4373.513639139139u,1.5 4373.514639139139u,0 4374.491179179179u,0 4374.492179179179u,1.5 4376.44625925926u,1.5 4376.44725925926u,0 4377.423799299299u,0 4377.4247992993u,1.5 4379.378879379379u,1.5 4379.379879379379u,0 4390.13181981982u,0 4390.13281981982u,1.5 4391.10935985986u,1.5 4391.11035985986u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.99706006006u,0 4395.99806006006u,1.5 4411.6377007007u,1.5 4411.638700700701u,0 4412.61524074074u,0 4412.61624074074u,1.5 4414.570320820821u,1.5 4414.571320820821u,0 4416.5254009009u,0 4416.526400900901u,1.5 4417.502940940941u,1.5 4417.503940940941u,0 4418.480480980981u,0 4418.481480980981u,1.5 4419.458021021021u,1.5 4419.459021021021u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4438.031281781782u,0 4438.032281781782u,1.5 4440.963901901901u,1.5 4440.964901901902u,0 4441.941441941942u,0 4441.942441941942u,1.5 4456.604542542542u,1.5 4456.605542542542u,0 4457.582082582582u,0 4457.583082582582u,1.5 4462.469782782783u,1.5 4462.470782782783u,0 4463.447322822823u,0 4463.448322822823u,1.5 4465.402402902902u,1.5 4465.403402902903u,0 4466.379942942943u,0 4466.380942942943u,1.5 4467.357482982983u,1.5 4467.358482982983u,0 4468.335023023023u,0 4468.336023023023u,1.5 4469.312563063063u,1.5 4469.313563063063u,0 4470.290103103103u,0 4470.2911031031035u,1.5 4471.267643143143u,1.5 4471.268643143143u,0 4472.245183183183u,0 4472.246183183183u,1.5 4473.222723223223u,1.5 4473.223723223223u,0 4476.155343343343u,0 4476.156343343343u,1.5 4478.1104234234235u,1.5 4478.111423423424u,0 4479.087963463464u,0 4479.088963463464u,1.5 4480.065503503503u,1.5 4480.066503503504u,0 4488.863363863864u,0 4488.864363863864u,1.5 4489.840903903903u,1.5 4489.841903903904u,0 4490.818443943944u,0 4490.819443943944u,1.5 4491.795983983984u,1.5 4491.796983983984u,0 4492.773524024024u,0 4492.774524024024u,1.5 4493.751064064064u,1.5 4493.752064064064u,0 4494.728604104104u,0 4494.7296041041045u,1.5 4495.706144144144u,1.5 4495.707144144144u,0 4502.5489244244245u,0 4502.549924424425u,1.5 4503.526464464465u,1.5 4503.527464464465u,0 4505.481544544544u,0 4505.482544544544u,1.5 4506.459084584585u,1.5 4506.460084584585u,0 4516.234484984985u,0 4516.235484984985u,1.5 4517.212025025025u,1.5 4517.213025025025u,0 4519.167105105105u,0 4519.1681051051055u,1.5 4520.144645145145u,1.5 4520.145645145145u,0 4521.122185185185u,0 4521.123185185185u,1.5 4523.077265265266u,1.5 4523.078265265266u,0 4524.054805305305u,0 4524.0558053053055u,1.5 4525.032345345345u,1.5 4525.033345345345u,0 4526.009885385385u,0 4526.010885385385u,1.5 4526.9874254254255u,1.5 4526.988425425426u,0 4528.942505505505u,0 4528.9435055055055u,1.5 4530.897585585586u,1.5 4530.898585585586u,0 4532.852665665666u,0 4532.853665665666u,1.5 4534.807745745745u,1.5 4534.808745745745u,0 4535.785285785786u,0 4535.786285785786u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4566.0890270270265u,0 4566.090027027027u,1.5 4567.066567067067u,1.5 4567.067567067067u,0 4584.662287787788u,0 4584.663287787788u,1.5 4585.6398278278275u,1.5 4585.640827827828u,0 4586.617367867868u,0 4586.618367867868u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4609.100788788789u,0 4609.101788788789u,1.5 4610.0783288288285u,1.5 4610.079328828829u,0 4620.83126926927u,0 4620.83226926927u,1.5 4623.763889389389u,1.5 4623.764889389389u,0 4624.741429429429u,0 4624.74242942943u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4636.471909909909u,0 4636.4729099099095u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4648.20239039039u,0 4648.20339039039u,1.5 4649.17993043043u,1.5 4649.180930430431u,0 4651.13501051051u,0 4651.1360105105105u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4675.573511511511u,0 4675.574511511511u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4696.101852352352u,0 4696.102852352352u,1.5 4698.056932432432u,1.5 4698.057932432433u,0 4699.034472472473u,0 4699.035472472473u,1.5 4700.989552552552u,1.5 4700.990552552552u,0 4701.967092592593u,0 4701.968092592593u,1.5 4704.899712712712u,1.5 4704.900712712712u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4715.652653153153u,0 4715.653653153153u,1.5 4716.630193193193u,1.5 4716.631193193193u,0 4718.585273273274u,0 4718.586273273274u,1.5 4719.562813313313u,1.5 4719.563813313313u,0 4720.540353353353u,0 4720.541353353353u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4731.293293793794u,0 4731.294293793794u,1.5 4732.270833833833u,1.5 4732.271833833834u,0 4739.113614114114u,0 4739.114614114114u,1.5 4740.091154154154u,1.5 4740.092154154154u,0 4741.068694194194u,0 4741.069694194194u,1.5 4742.046234234233u,1.5 4742.047234234234u,0 4743.023774274275u,0 4743.024774274275u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4759.6419549549555u,0 4759.642954954956u,1.5 4760.619494994995u,1.5 4760.620494994995u,0 4761.597035035034u,0 4761.598035035035u,1.5 4768.439815315315u,1.5 4768.440815315315u,0 4769.4173553553555u,0 4769.418355355356u,1.5 4771.372435435435u,1.5 4771.373435435436u,0 4782.125375875876u,0 4782.126375875876u,1.5 4783.102915915916u,1.5 4783.103915915916u,0 4784.0804559559565u,0 4784.081455955957u,1.5 4793.8558563563565u,1.5 4793.856856356357u,0 4802.653716716716u,0 4802.654716716716u,1.5 4803.6312567567575u,1.5 4803.632256756758u,0 4805.586336836836u,0 4805.587336836837u,1.5 4806.563876876877u,1.5 4806.564876876877u,0 4807.541416916917u,0 4807.542416916917u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4825.137137637637u,0 4825.138137637638u,1.5 4826.114677677678u,1.5 4826.115677677678u,0 4828.069757757758u,0 4828.070757757759u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4840.777778278279u,0 4840.778778278279u,1.5 4841.755318318318u,1.5 4841.756318318318u,0 4848.598098598599u,0 4848.599098598599u,1.5 4849.575638638638u,1.5 4849.5766386386385u,0 4852.508258758759u,0 4852.50925875876u,1.5 4863.261199199199u,1.5 4863.262199199199u,0 4864.238739239238u,0 4864.239739239239u,1.5 4866.193819319319u,1.5 4866.194819319319u,0 4875.969219719719u,0 4875.970219719719u,1.5 4876.94675975976u,1.5 4876.947759759761u,0 4877.9242997998u,0 4877.9252997998u,1.5 4878.901839839839u,1.5 4878.9028398398395u,0 4879.87937987988u,0 4879.88037987988u,1.5 4880.85691991992u,1.5 4880.85791991992u,0 4881.83445995996u,0 4881.835459959961u,1.5 4891.6098603603605u,1.5 4891.610860360361u,0 4892.5874004004u,0 4892.5884004004u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4894.542480480481u,0 4894.543480480481u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4898.45264064064u,0 4898.4536406406405u,1.5 4899.430180680681u,1.5 4899.431180680681u,0 4912.138201201201u,0 4912.139201201201u,1.5 4913.11574124124u,1.5 4913.116741241241u,0 4914.093281281282u,0 4914.094281281282u,1.5 4915.070821321321u,1.5 4915.071821321321u,0 4916.0483613613615u,0 4916.049361361362u,1.5 4917.025901401401u,1.5 4917.026901401401u,0 4918.003441441441u,0 4918.0044414414415u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4938.531782282283u,1.5 4938.532782282283u,0 4940.486862362362u,0 4940.487862362363u,1.5 4941.464402402402u,1.5 4941.465402402402u,0 4965.902903403403u,0 4965.903903403403u,1.5 4966.880443443443u,1.5 4966.8814434434435u,0 4968.835523523523u,0 4968.836523523523u,1.5 4970.790603603604u,1.5 4970.791603603604u,0 4971.768143643643u,0 4971.7691436436435u,1.5 4972.745683683684u,1.5 4972.746683683684u,0 4973.723223723723u,0 4973.724223723723u,1.5 4974.700763763764u,1.5 4974.701763763765u,0 4975.678303803804u,0 4975.679303803804u,1.5 4976.655843843843u,1.5 4976.6568438438435u,0 4977.633383883884u,0 4977.634383883884u,1.5 4979.588463963964u,1.5 4979.589463963965u,0 4980.566004004004u,0 4980.567004004004u,1.5 4983.498624124124u,1.5 4983.499624124124u,0 4984.476164164164u,0 4984.477164164165u,1.5 4986.431244244243u,1.5 4986.4322442442435u,0 4987.408784284285u,0 4987.409784284285u,1.5 4989.363864364364u,1.5 4989.364864364365u,0 4990.341404404404u,0 4990.342404404404u,1.5 4992.296484484485u,1.5 4992.297484484485u,0 4993.274024524524u,0 4993.275024524524u,1.5 4996.206644644644u,1.5 4996.2076446446445u,0 4997.184184684685u,0 4997.185184684685u,1.5 5007.937125125125u,1.5 5007.938125125125u,0 5008.914665165165u,0 5008.915665165166u,1.5 5014.779905405405u,1.5 5014.780905405405u,0 5015.757445445445u,0 5015.758445445445u,1.5 5016.734985485486u,1.5 5016.735985485486u,0 5017.712525525525u,0 5017.713525525525u,1.5 5021.622685685686u,1.5 5021.623685685686u,0 5022.600225725725u,0 5022.601225725725u,1.5 5024.555305805806u,1.5 5024.556305805806u,0 5025.532845845845u,0 5025.5338458458455u,1.5 5027.487925925926u,1.5 5027.488925925926u,0 5028.465465965966u,0 5028.466465965967u,1.5 5029.443006006006u,1.5 5029.444006006006u,0 5030.420546046045u,0 5030.4215460460455u,1.5 5031.398086086087u,1.5 5031.399086086087u,0 5033.353166166166u,0 5033.354166166167u,1.5 5035.308246246245u,1.5 5035.3092462462455u,0 5057.791667167167u,0 5057.792667167168u,1.5 5058.769207207207u,1.5 5058.770207207207u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5064.634447447447u,0 5064.635447447447u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5086.140328328328u,1.5 5086.141328328328u,0 5087.117868368368u,0 5087.118868368369u,1.5 5088.095408408408u,1.5 5088.096408408408u,0 5090.050488488489u,0 5090.051488488489u,1.5 5092.005568568568u,1.5 5092.006568568569u,0 5092.983108608609u,0 5092.984108608609u,1.5 5093.960648648648u,1.5 5093.961648648648u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5120.354229729729u,1.5 5120.355229729729u,0 5121.33176976977u,0 5121.3327697697705u,1.5 5123.286849849849u,1.5 5123.287849849849u,0 5124.26438988989u,0 5124.26538988989u,1.5 5125.24192992993u,1.5 5125.24292992993u,0 5135.01733033033u,0 5135.01833033033u,1.5 5135.99487037037u,1.5 5135.9958703703705u,0 5136.97241041041u,0 5136.97341041041u,1.5 5149.680430930931u,1.5 5149.681430930931u,0 5150.657970970971u,0 5150.6589709709715u,1.5 5152.61305105105u,1.5 5152.61405105105u,0 5160.433371371371u,0 5160.4343713713715u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5162.388451451451u,0 5162.389451451451u,1.5 5171.186311811812u,1.5 5171.187311811812u,0 5172.163851851851u,0 5172.164851851851u,1.5 5174.118931931932u,1.5 5174.119931931932u,0 5176.074012012012u,0 5176.075012012012u,1.5 5177.051552052051u,1.5 5177.052552052051u,0 5186.826952452452u,0 5186.827952452452u,1.5 5194.647272772773u,1.5 5194.648272772773u,0 5195.624812812813u,0 5195.625812812813u,1.5 5198.557432932933u,1.5 5198.558432932933u,0 5208.332833333333u,0 5208.333833333333u,1.5 5218.108233733733u,1.5 5218.109233733733u,0 5220.063313813814u,0 5220.064313813814u,1.5 5221.040853853853u,1.5 5221.041853853853u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5232.771334334334u,0 5232.772334334334u,1.5 5237.659034534534u,1.5 5237.660034534534u,0 5238.636574574574u,0 5238.6375745745745u,1.5 5240.591654654654u,1.5 5240.592654654654u,0 5250.367055055054u,0 5250.368055055054u,1.5 5258.187375375375u,1.5 5258.1883753753755u,0 5259.164915415415u,0 5259.165915415415u,1.5 5260.142455455456u,1.5 5260.143455455456u,0 5261.1199954954955u,0 5261.120995495496u,1.5 5262.097535535535u,1.5 5262.098535535535u,0 5271.872935935936u,0 5271.873935935936u,1.5 5280.670796296296u,1.5 5280.671796296297u,0 5281.648336336336u,0 5281.649336336336u,1.5 5282.625876376376u,1.5 5282.6268763763765u,0 5283.603416416417u,0 5283.604416416417u,1.5 5284.580956456457u,1.5 5284.581956456457u,0 5289.468656656657u,0 5289.469656656657u,1.5 5290.4461966966965u,1.5 5290.447196696697u,0 5292.401276776777u,0 5292.402276776777u,1.5 5294.356356856857u,1.5 5294.357356856857u,0 5295.3338968968965u,0 5295.334896896897u,1.5 5299.244057057057u,1.5 5299.245057057057u,0 5300.221597097097u,0 5300.222597097098u,1.5 5302.176677177177u,1.5 5302.177677177177u,0 5303.154217217217u,0 5303.155217217217u,1.5 5304.131757257258u,1.5 5304.132757257258u,0 5305.109297297297u,0 5305.110297297298u,1.5 5306.086837337337u,1.5 5306.087837337337u,0 5312.929617617618u,0 5312.930617617618u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5326.615178178178u,1.5 5326.616178178178u,0 5327.592718218218u,0 5327.593718218218u,1.5 5328.570258258259u,1.5 5328.571258258259u,0 5337.368118618619u,0 5337.369118618619u,1.5 5338.345658658659u,1.5 5338.346658658659u,0 5339.323198698698u,0 5339.324198698699u,1.5 5351.053679179179u,1.5 5351.054679179179u,0 5352.031219219219u,0 5352.032219219219u,1.5 5353.00875925926u,1.5 5353.00975925926u,0 5354.963839339339u,0 5354.964839339339u,1.5 5355.941379379379u,1.5 5355.942379379379u,0 5362.78415965966u,0 5362.78515965966u,1.5 5363.761699699699u,1.5 5363.7626996997u,0 5364.739239739739u,0 5364.740239739739u,1.5 5366.69431981982u,1.5 5366.69531981982u,0 5367.67185985986u,0 5367.67285985986u,1.5 5376.46972022022u,1.5 5376.47072022022u,0 5377.447260260261u,0 5377.448260260261u,1.5 5378.4248003003u,1.5 5378.425800300301u,0 5394.065440940941u,0 5394.066440940941u,1.5 5395.042980980981u,1.5 5395.043980980981u,0 5396.020521021021u,0 5396.021521021021u,1.5 5396.998061061061u,1.5 5396.999061061061u,0 5397.975601101101u,0 5397.976601101102u,1.5 5398.953141141141u,1.5 5398.954141141141u,0 5399.930681181181u,0 5399.931681181181u,1.5 5407.751001501501u,1.5 5407.752001501502u,0 5408.728541541541u,0 5408.729541541541u,1.5 5410.683621621622u,1.5 5410.684621621622u,0 5411.661161661662u,0 5411.662161661662u,1.5 5413.616241741741u,1.5 5413.617241741741u,0 5430.2344224224225u,0 5430.235422422423u,1.5 5431.211962462463u,1.5 5431.212962462463u,0 5432.189502502502u,0 5432.190502502503u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5438.054742742742u,1.5 5438.055742742742u,0 5439.032282782783u,0 5439.033282782783u,1.5 5440.009822822823u,1.5 5440.010822822823u,0 5440.987362862863u,0 5440.988362862863u,1.5 5444.897523023023u,1.5 5444.898523023023u,0 5445.875063063063u,0 5445.876063063063u,1.5 5461.515703703703u,1.5 5461.516703703704u,0 5462.493243743743u,0 5462.494243743743u,1.5 5464.448323823824u,1.5 5464.449323823824u,0 5465.425863863864u,0 5465.426863863864u,1.5 5470.313564064064u,1.5 5470.314564064064u,0 5471.291104104104u,0 5471.2921041041045u,1.5 5473.246184184184u,1.5 5473.247184184184u,0 5474.223724224224u,0 5474.224724224224u,1.5 5475.201264264265u,1.5 5475.202264264265u,0 5478.133884384384u,0 5478.134884384384u,1.5 5479.1114244244245u,1.5 5479.112424424425u,0 5481.066504504504u,0 5481.0675045045045u,1.5 5482.044044544544u,1.5 5482.045044544544u,0 5483.021584584585u,0 5483.022584584585u,1.5 5483.9991246246245u,1.5 5484.000124624625u,0 5484.976664664665u,0 5484.977664664665u,1.5 5485.954204704704u,1.5 5485.955204704705u,0 5488.8868248248245u,0 5488.887824824825u,1.5 5489.864364864865u,1.5 5489.865364864865u,0 5492.796984984985u,0 5492.797984984985u,1.5 5493.774525025025u,1.5 5493.775525025025u,0 5495.729605105105u,0 5495.7306051051055u,1.5 5496.707145145145u,1.5 5496.708145145145u,0 5499.639765265266u,0 5499.640765265266u,1.5 5500.617305305305u,1.5 5500.6183053053055u,0 5510.392705705705u,0 5510.3937057057055u,1.5 5511.370245745745u,1.5 5511.371245745745u,0 5515.280405905905u,0 5515.281405905906u,1.5 5516.257945945946u,1.5 5516.258945945946u,0 5517.235485985986u,0 5517.236485985986u,1.5 5518.213026026026u,1.5 5518.214026026026u,0 5520.168106106106u,0 5520.1691061061065u,1.5 5521.145646146146u,1.5 5521.146646146146u,0 5524.078266266267u,0 5524.079266266267u,1.5 5525.055806306306u,1.5 5525.0568063063065u,0 5526.033346346346u,0 5526.034346346346u,1.5 5527.010886386386u,1.5 5527.011886386386u,0 5527.9884264264265u,0 5527.989426426427u,1.5 5529.943506506506u,1.5 5529.9445065065065u,0 5530.921046546546u,0 5530.922046546546u,1.5 5531.898586586587u,1.5 5531.899586586587u,0 5533.853666666667u,0 5533.854666666667u,1.5 5540.696446946947u,1.5 5540.697446946947u,0 5541.673986986987u,0 5541.674986986987u,1.5 5558.292167667668u,1.5 5558.293167667668u,0 5559.269707707707u,0 5559.2707077077075u,1.5 5562.2023278278275u,1.5 5562.203327827828u,0 5563.179867867868u,0 5563.180867867868u,1.5 5566.112487987988u,1.5 5566.113487987988u,0 5567.0900280280275u,0 5567.091028028028u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5570.022648148148u,0 5570.023648148148u,1.5 5571.000188188188u,1.5 5571.001188188188u,0 5584.685748748749u,0 5584.686748748749u,1.5 5585.663288788789u,1.5 5585.664288788789u,0 5586.6408288288285u,0 5586.641828828829u,1.5 5587.618368868869u,1.5 5587.619368868869u,0 5589.573448948949u,0 5589.574448948949u,1.5 5600.326389389389u,1.5 5600.327389389389u,0 5601.303929429429u,0 5601.30492942943u,1.5 5605.21408958959u,1.5 5605.21508958959u,0 5608.146709709709u,0 5608.1477097097095u,1.5 5609.12424974975u,1.5 5609.12524974975u,0 5620.8547302302295u,0 5620.85573023023u,1.5 5621.832270270271u,1.5 5621.833270270271u,0 5623.78735035035u,0 5623.78835035035u,1.5 5633.562750750751u,1.5 5633.563750750751u,0 5634.540290790791u,0 5634.541290790791u,1.5 5636.495370870871u,1.5 5636.496370870871u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5638.450450950951u,1.5 5638.451450950951u,0 5648.225851351351u,0 5648.226851351351u,1.5 5649.203391391391u,1.5 5649.204391391391u,0 5650.180931431431u,0 5650.181931431432u,1.5 5651.158471471472u,1.5 5651.159471471472u,0 5652.136011511511u,0 5652.137011511511u,1.5 5653.113551551551u,1.5 5653.114551551551u,0 5654.091091591592u,0 5654.092091591592u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5664.8440320320315u,0 5664.845032032032u,1.5 5665.821572072072u,1.5 5665.822572072072u,0 5675.596972472473u,0 5675.597972472473u,1.5 5676.574512512512u,1.5 5676.575512512512u,0 5677.552052552552u,0 5677.553052552552u,1.5 5682.439752752753u,1.5 5682.440752752753u,0 5683.417292792793u,0 5683.418292792793u,1.5 5685.372372872873u,1.5 5685.373372872873u,0 5688.304992992993u,0 5688.305992992993u,1.5 5689.282533033032u,1.5 5689.283533033033u,0 5695.147773273274u,0 5695.148773273274u,1.5 5696.125313313313u,1.5 5696.126313313313u,0 5699.057933433433u,0 5699.058933433434u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5715.676114114114u,0 5715.677114114114u,1.5 5716.653654154154u,1.5 5716.654654154154u,0 5718.608734234233u,0 5718.609734234234u,1.5 5727.406594594595u,1.5 5727.407594594595u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5740.114615115115u,0 5740.115615115115u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 5758.687875875876u,0 5758.688875875876u,1.5 5759.665415915916u,1.5 5759.666415915916u,0 5760.6429559559565u,0 5760.643955955957u,1.5 5761.620495995996u,1.5 5761.621495995996u,0 5762.598036036035u,0 5762.599036036036u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5772.373436436436u,1.5 5772.374436436437u,0 5778.238676676677u,0 5778.239676676677u,1.5 5779.216216716716u,1.5 5779.217216716716u,0 5781.171296796797u,0 5781.172296796797u,1.5 5782.148836836836u,1.5 5782.149836836837u,0 5783.126376876877u,0 5783.127376876877u,1.5 5788.991617117117u,1.5 5788.992617117117u,0 5789.9691571571575u,0 5789.970157157158u,1.5 5790.946697197197u,1.5 5790.947697197197u,0 5792.901777277278u,0 5792.902777277278u,1.5 5793.879317317317u,1.5 5793.880317317317u,0 5800.722097597598u,0 5800.723097597598u,1.5 5801.699637637637u,1.5 5801.700637637638u,0 5802.677177677678u,0 5802.678177677678u,1.5 5813.430118118118u,1.5 5813.431118118118u,0 5815.385198198198u,0 5815.386198198198u,1.5 5816.362738238237u,1.5 5816.363738238238u,0 5825.160598598599u,0 5825.161598598599u,1.5 5827.115678678679u,1.5 5827.116678678679u,0 5829.070758758759u,0 5829.07175875876u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5838.8461591591595u,0 5838.84715915916u,1.5 5840.801239239238u,1.5 5840.802239239239u,0 5849.5990995996u,0 5849.6000995996u,1.5 5851.55417967968u,1.5 5851.55517967968u,0 5852.531719719719u,0 5852.532719719719u,1.5 5859.3745u,1.5 5859.3755u,0 5860.352040040039u,0 5860.35304004004u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5863.2846601601605u,0 5863.285660160161u,1.5 5864.2622002002u,1.5 5864.2632002002u,0 5876.97022072072u,0 5876.97122072072u,1.5 5877.947760760761u,1.5 5877.948760760762u,0 5878.925300800801u,0 5878.926300800801u,1.5 5880.880380880881u,1.5 5880.881380880881u,0 5882.835460960961u,0 5882.836460960962u,1.5 5888.700701201201u,1.5 5888.701701201201u,0 5889.67824124124u,0 5889.679241241241u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5899.453641641641u,0 5899.4546416416415u,1.5 5900.431181681682u,1.5 5900.432181681682u,0 5908.251502002002u,0 5908.252502002002u,1.5 5909.229042042041u,1.5 5909.2300420420415u,0 5910.206582082082u,0 5910.207582082082u,1.5 5911.184122122122u,1.5 5911.185122122122u,0 5912.161662162162u,0 5912.162662162163u,1.5 5932.690003003003u,1.5 5932.691003003003u,0 5933.667543043042u,0 5933.6685430430425u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5936.600163163163u,0 5936.601163163164u,1.5 5938.555243243242u,1.5 5938.5562432432425u,0 5958.106044044043u,0 5958.1070440440435u,1.5 5959.083584084084u,1.5 5959.084584084084u,0 5960.061124124124u,0 5960.062124124124u,1.5 5961.038664164164u,1.5 5961.039664164165u,0 5963.971284284285u,0 5963.972284284285u,1.5 5964.948824324324u,1.5 5964.949824324324u,0 5968.858984484485u,0 5968.859984484485u,1.5 5970.814064564564u,1.5 5970.815064564565u,0 5971.791604604605u,0 5971.792604604605u,1.5 5972.769144644644u,1.5 5972.7701446446445u,0 5973.746684684685u,0 5973.747684684685u,1.5 5979.611924924925u,1.5 5979.612924924925u,0 5980.589464964965u,0 5980.590464964966u,1.5 5983.522085085086u,1.5 5983.523085085086u,0 5984.499625125125u,0 5984.500625125125u,1.5 6006.005506006006u,1.5 6006.006506006006u,0 6006.983046046045u,0 6006.9840460460455u,1.5 6012.848286286287u,1.5 6012.849286286287u,0 6013.825826326326u,0 6013.826826326326u,1.5 6017.735986486487u,1.5 6017.736986486487u,0 6018.713526526526u,0 6018.714526526526u,1.5 6023.601226726726u,1.5 6023.602226726726u,0 6024.578766766767u,0 6024.5797667667675u,1.5 6028.488926926927u,1.5 6028.489926926927u,0 6029.466466966967u,0 6029.467466966968u,1.5 6030.444007007007u,1.5 6030.445007007007u,0 6032.3990870870875u,0 6032.400087087088u,1.5 6033.376627127127u,1.5 6033.377627127127u,0 6036.309247247247u,0 6036.310247247247u,1.5 6037.286787287288u,1.5 6037.287787287288u,0 6055.860048048047u,0 6055.861048048047u,1.5 6056.8375880880885u,1.5 6056.838588088089u,0 6059.770208208208u,0 6059.771208208208u,1.5 6060.747748248248u,1.5 6060.748748248248u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6068.568068568568u,1.5 6068.569068568569u,0 6070.523148648648u,0 6070.524148648648u,1.5 6071.500688688689u,1.5 6071.501688688689u,0 6072.478228728728u,0 6072.479228728728u,1.5 6074.433308808809u,1.5 6074.434308808809u,0 6075.410848848848u,0 6075.411848848848u,1.5 6087.141329329329u,1.5 6087.142329329329u,0 6088.118869369369u,0 6088.11986936937u,1.5 6090.073949449449u,1.5 6090.074949449449u,0 6101.80442992993u,0 6101.80542992993u,1.5 6102.78196996997u,1.5 6102.7829699699705u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6106.69213013013u,0 6106.69313013013u,1.5 6107.66967017017u,1.5 6107.6706701701705u,0 6108.64721021021u,0 6108.64821021021u,1.5 6118.422610610611u,1.5 6118.423610610611u,0 6119.40015065065u,0 6119.40115065065u,1.5 6120.3776906906905u,1.5 6120.378690690691u,0 6136.018331331331u,0 6136.019331331331u,1.5 6137.973411411411u,1.5 6137.974411411411u,0 6138.950951451451u,0 6138.951951451451u,1.5 6139.9284914914915u,1.5 6139.929491491492u,0 6140.906031531531u,0 6140.907031531531u,1.5 6147.748811811812u,1.5 6147.749811811812u,0 6148.726351851851u,0 6148.727351851851u,1.5 6151.658971971972u,1.5 6151.6599719719725u,0 6152.636512012012u,0 6152.637512012012u,1.5 6153.614052052051u,1.5 6153.615052052051u,0 6159.4792922922925u,0 6159.480292292293u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6162.411912412412u,0 6162.412912412412u,1.5 6172.187312812813u,1.5 6172.188312812813u,0 6173.164852852852u,0 6173.165852852852u,1.5 6175.119932932933u,1.5 6175.120932932933u,0 6176.097472972973u,0 6176.0984729729735u,1.5 6177.075013013013u,1.5 6177.076013013013u,0 6184.895333333333u,0 6184.896333333333u,1.5 6185.872873373373u,1.5 6185.8738733733735u,0 6186.850413413413u,0 6186.851413413413u,1.5 6197.603353853853u,1.5 6197.604353853853u,0 6200.535973973974u,0 6200.536973973974u,1.5 6201.513514014014u,1.5 6201.514514014014u,0 6208.3562942942945u,0 6208.357294294295u,1.5 6215.199074574574u,1.5 6215.2000745745745u,0 6216.176614614615u,0 6216.177614614615u,1.5 6219.109234734734u,1.5 6219.110234734734u,0 6220.086774774775u,0 6220.087774774775u,1.5 6221.064314814815u,1.5 6221.065314814815u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6232.794795295295u,0 6232.795795295296u,1.5 6239.637575575575u,1.5 6239.6385755755755u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6256.255756256256u,1.5 6256.256756256256u,0 6257.233296296296u,0 6257.234296296297u,1.5 6260.165916416417u,1.5 6260.166916416417u,0 6261.143456456457u,0 6261.144456456457u,1.5 6262.120996496496u,1.5 6262.121996496497u,0 6268.963776776777u,0 6268.964776776777u,1.5 6269.941316816817u,1.5 6269.942316816817u,0 6270.918856856857u,0 6270.919856856857u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6272.873936936937u,0 6272.874936936937u,1.5 6278.739177177177u,1.5 6278.740177177177u,0 6279.716717217217u,0 6279.717717217217u,1.5 6282.649337337337u,1.5 6282.650337337337u,0 6283.626877377377u,0 6283.627877377377u,1.5 6284.604417417418u,1.5 6284.605417417418u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6291.447197697697u,0 6291.448197697698u,1.5 6304.155218218218u,1.5 6304.156218218218u,0 6305.132758258259u,0 6305.133758258259u,1.5 6306.110298298298u,1.5 6306.111298298299u,0 6307.087838338338u,0 6307.088838338338u,1.5 6308.065378378378u,1.5 6308.066378378378u,0 6313.930618618619u,0 6313.931618618619u,1.5 6314.908158658659u,1.5 6314.909158658659u,0 6315.885698698698u,0 6315.886698698699u,1.5 6317.840778778779u,1.5 6317.841778778779u,0 6318.818318818819u,0 6318.819318818819u,1.5 6326.638639139139u,1.5 6326.639639139139u,0 6337.391579579579u,0 6337.392579579579u,1.5 6339.34665965966u,1.5 6339.34765965966u,0 6340.324199699699u,0 6340.3251996997u,1.5 6342.27927977978u,1.5 6342.28027977978u,0 6343.25681981982u,0 6343.25781981982u,1.5 6350.0996001001u,1.5 6350.100600100101u,0 6351.07714014014u,0 6351.07814014014u,1.5 6352.05468018018u,1.5 6352.05568018018u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6363.785160660661u,0 6363.786160660661u,1.5 6379.425801301301u,1.5 6379.426801301302u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6397.021522022022u,0 6397.022522022022u,1.5 6406.7969224224225u,1.5 6406.797922422423u,0 6407.774462462463u,0 6407.775462462463u,1.5 6410.707082582582u,1.5 6410.708082582582u,0 6411.684622622623u,0 6411.685622622623u,1.5 6414.617242742742u,1.5 6414.618242742742u,0 6416.572322822823u,0 6416.573322822823u,1.5 6417.549862862863u,1.5 6417.550862862863u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6437.100663663664u,0 6437.101663663664u,1.5 6446.876064064064u,1.5 6446.877064064064u,0 6447.853604104104u,0 6447.8546041041045u,1.5 6463.494244744744u,1.5 6463.495244744744u,0 6464.471784784785u,0 6464.472784784785u,1.5 6465.4493248248245u,1.5 6465.450324824825u,0 6466.426864864865u,0 6466.427864864865u,1.5 6468.381944944945u,1.5 6468.382944944945u,0 6469.359484984985u,0 6469.360484984985u,1.5 6471.314565065065u,1.5 6471.315565065065u,0 6472.292105105105u,0 6472.2931051051055u,1.5 6474.247185185185u,1.5 6474.248185185185u,0 6476.202265265266u,0 6476.203265265266u,1.5 6477.179805305305u,1.5 6477.1808053053055u,0 6484.022585585586u,0 6484.023585585586u,1.5 6485.0001256256255u,1.5 6485.001125625626u,0 6488.910285785786u,0 6488.911285785786u,1.5 6489.8878258258255u,1.5 6489.888825825826u,0 6500.640766266267u,0 6500.641766266267u,1.5 6501.618306306306u,1.5 6501.6193063063065u,0 6511.393706706706u,0 6511.3947067067065u,1.5 6512.371246746747u,1.5 6512.372246746747u,0 6517.258946946947u,0 6517.259946946947u,1.5 6518.236486986987u,1.5 6518.237486986987u,0 6520.191567067067u,0 6520.192567067067u,1.5 6521.169107107107u,1.5 6521.1701071071075u,0 6525.079267267268u,0 6525.080267267268u,1.5 6527.034347347347u,1.5 6527.035347347347u,0 6528.9894274274275u,0 6528.990427427428u,1.5 6532.899587587588u,1.5 6532.900587587588u,0 6533.8771276276275u,0 6533.878127627628u,1.5 6535.832207707707u,1.5 6535.8332077077075u,0 6536.809747747748u,0 6536.810747747748u,1.5 6562.225788788789u,1.5 6562.226788788789u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6565.158408908908u,0 6565.1594089089085u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6568.0910290290285u,0 6568.092029029029u,1.5 6569.068569069069u,1.5 6569.069569069069u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.001189189189u,1.5 6572.002189189189u,0 6586.66428978979u,0 6586.66528978979u,1.5 6587.6418298298295u,1.5 6587.64282982983u,0 6588.61936986987u,0 6588.62036986987u,1.5 6590.57444994995u,1.5 6590.57544994995u,0 6591.55198998999u,0 6591.55298998999u,1.5 6600.34985035035u,1.5 6600.35085035035u,0 6601.32739039039u,0 6601.32839039039u,1.5 6604.26001051051u,1.5 6604.2610105105105u,0 6606.215090590591u,0 6606.216090590591u,1.5 6607.19263063063u,1.5 6607.193630630631u,0 6618.923111111111u,0 6618.924111111111u,1.5 6619.900651151151u,1.5 6619.901651151151u,0 6621.8557312312305u,0 6621.856731231231u,1.5 6623.810811311311u,1.5 6623.811811311311u,0 6624.788351351351u,0 6624.789351351351u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6637.496371871872u,1.5 6637.497371871872u,0 6638.473911911911u,0 6638.4749119119115u,1.5 6639.451451951952u,1.5 6639.452451951952u,0 6649.226852352352u,0 6649.227852352352u,1.5 6650.204392392392u,1.5 6650.205392392392u,0 6651.181932432432u,0 6651.182932432433u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6664.867492992993u,0 6664.868492992993u,1.5 6665.845033033032u,1.5 6665.846033033033u,0 6672.687813313313u,0 6672.688813313313u,1.5 6673.665353353353u,1.5 6673.666353353353u,0 6674.642893393393u,0 6674.643893393393u,1.5 6676.597973473474u,1.5 6676.598973473474u,0 6677.575513513513u,0 6677.576513513513u,1.5 6685.395833833833u,1.5 6685.396833833834u,0 6693.216154154154u,0 6693.217154154154u,1.5 6694.193694194194u,1.5 6694.194694194194u,0 6698.103854354354u,0 6698.104854354354u,1.5 6705.924174674675u,1.5 6705.925174674675u,0 6706.901714714714u,0 6706.902714714714u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6708.856794794795u,0 6708.857794794795u,1.5 6709.834334834834u,1.5 6709.835334834835u,0 6718.632195195195u,0 6718.633195195195u,1.5 6719.609735235234u,1.5 6719.610735235235u,0 6720.587275275276u,0 6720.588275275276u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6727.430055555555u,0 6727.431055555555u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6741.115616116116u,0 6741.116616116116u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6752.846096596597u,1.5 6752.847096596597u,0 6761.6439569569575u,0 6761.644956956958u,1.5 6768.486737237236u,1.5 6768.487737237237u,0 6769.464277277278u,0 6769.465277277278u,1.5 6771.4193573573575u,1.5 6771.420357357358u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6780.217217717717u,0 6780.218217717717u,1.5 6782.172297797798u,1.5 6782.173297797798u,0 6783.149837837837u,0 6783.150837837838u,1.5 6791.947698198198u,1.5 6791.948698198198u,0 6802.700638638638u,0 6802.7016386386385u,1.5 6803.678178678679u,1.5 6803.679178678679u,0 6804.655718718718u,0 6804.656718718718u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6814.431119119119u,0 6814.432119119119u,1.5 6815.4086591591595u,1.5 6815.40965915916u,0 6823.22897947948u,0 6823.22997947948u,1.5 6824.206519519519u,1.5 6824.207519519519u,0 6826.1615995996u,0 6826.1625995996u,1.5 6827.139139639639u,1.5 6827.1401396396395u,0 6828.11667967968u,0 6828.11767967968u,1.5 6835.937u,1.5 6835.938u,0 6837.89208008008u,0 6837.89308008008u,1.5 6839.8471601601605u,1.5 6839.848160160161u,0 6848.64502052052u,0 6848.64602052052u,1.5 6849.6225605605605u,1.5 6849.623560560561u,0 6851.57764064064u,0 6851.5786406406405u,1.5 6854.510260760761u,1.5 6854.511260760762u,0 6855.487800800801u,0 6855.488800800801u,1.5 6860.375501001001u,1.5 6860.376501001001u,0 6861.35304104104u,0 6861.354041041041u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6866.24074124124u,0 6866.241741241241u,1.5 6867.218281281282u,1.5 6867.219281281282u,0 6876.016141641641u,0 6876.0171416416415u,1.5 6876.993681681682u,1.5 6876.994681681682u,0 6878.948761761762u,0 6878.949761761763u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6893.611862362362u,0 6893.612862362363u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6908.274962962963u,0 6908.275962962964u,1.5 6909.252503003003u,1.5 6909.253503003003u,0 6912.185123123123u,0 6912.186123123123u,1.5 6913.162663163163u,1.5 6913.163663163164u,0 6914.140203203203u,0 6914.141203203203u,1.5 6932.713463963964u,1.5 6932.714463963965u,0 6933.691004004004u,0 6933.692004004004u,1.5 6934.668544044043u,1.5 6934.6695440440435u,0 6935.646084084084u,0 6935.647084084084u,1.5 6936.623624124124u,1.5 6936.624624124124u,0 6938.578704204204u,0 6938.579704204204u,1.5 6939.556244244243u,1.5 6939.5572442442435u,0 6942.488864364364u,0 6942.489864364365u,1.5 6943.466404404404u,1.5 6943.467404404404u,0 6962.039665165165u,0 6962.040665165166u,1.5 6963.017205205205u,1.5 6963.018205205205u,0 6963.994745245244u,0 6963.9957452452445u,1.5 6964.972285285286u,1.5 6964.973285285286u,0 6967.904905405405u,0 6967.905905405405u,1.5 6968.882445445445u,1.5 6968.883445445445u,0 6969.859985485486u,0 6969.860985485486u,1.5 6970.837525525525u,1.5 6970.838525525525u,0 6971.815065565565u,0 6971.816065565566u,1.5 6972.792605605606u,1.5 6972.793605605606u,0 6973.770145645645u,0 6973.771145645645u,1.5 6974.747685685686u,1.5 6974.748685685686u,0 6976.702765765766u,0 6976.703765765767u,1.5 6978.657845845845u,1.5 6978.6588458458455u,0 6979.635385885886u,0 6979.636385885886u,1.5 6981.590465965966u,1.5 6981.591465965967u,0 6982.568006006006u,0 6982.569006006006u,1.5 6986.478166166166u,1.5 6986.479166166167u,0 6987.455706206206u,0 6987.456706206206u,1.5 6989.410786286287u,1.5 6989.411786286287u,0 6990.388326326326u,0 6990.389326326326u,1.5 6991.365866366366u,1.5 6991.366866366367u,0 6992.343406406406u,0 6992.344406406406u,1.5 6994.298486486487u,1.5 6994.299486486487u,0 6995.276026526526u,0 6995.277026526526u,1.5
vbb13 bb13 0 pwl 0,1.5  58.6519024024024u,1.5 58.652902402402404u,0 59.62944244244244u,0 59.630442442442444u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 104.59628428428428u,0 104.59728428428429u,1.5 106.55136436436436u,1.5 106.55236436436437u,0 107.5289044044044u,0 107.5299044044044u,1.5 109.48398448448448u,1.5 109.48498448448449u,0 110.46152452452452u,0 110.46252452452453u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 136.85510560560562u,0 136.8561056056056u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 164.22622672672674u,0 164.2272267267267u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 185.73210760760762u,0 185.7331076076076u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 188.66472772772775u,1.5 188.66572772772773u,0 207.2379884884885u,0 207.23898848848847u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 210.17060860860863u,0 210.1716086086086u,1.5 229.72140940940943u,1.5 229.7224094094094u,0 230.69894944944946u,0 230.69994944944943u,1.5 231.6764894894895u,1.5 231.6774894894895u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 270.77809109109114u,1.5 270.7790910910911u,0 271.75563113113117u,0 271.75663113113114u,1.5 272.73317117117114u,1.5 272.7341711711711u,0 289.35135185185186u,0 289.35235185185184u,1.5 290.32889189189194u,1.5 290.3298918918919u,0 294.23905205205205u,0 294.240052052052u,1.5 313.78985285285285u,1.5 313.7908528528528u,0 314.76739289289293u,0 314.7683928928929u,1.5 315.74493293293295u,1.5 315.74593293293293u,0 317.700013013013u,0 317.701013013013u,1.5 318.67755305305303u,1.5 318.678553053053u,0 335.2957337337337u,0 335.2967337337337u,1.5 336.2732737737738u,1.5 336.27427377377376u,0 337.2508138138138u,0 337.2518138138138u,1.5 338.2283538538539u,1.5 338.22935385385387u,0 340.18343393393394u,0 340.1844339339339u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 389.06043593593597u,0 389.06143593593595u,1.5 390.037975975976u,1.5 390.038975975976u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 395.90321621621626u,0 395.90421621621624u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 432.07219769769773u,1.5 432.0731976976977u,0 433.04973773773776u,0 433.05073773773773u,1.5 434.0272777777778u,1.5 434.02827777777776u,0 435.00481781781787u,0 435.00581781781784u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 437.93743793793794u,0 437.9384379379379u,1.5 438.91497797797797u,1.5 438.91597797797795u,0 560.1299429429429u,0 560.1309429429429u,1.5 561.107482982983u,1.5 561.108482982983u,0 563.0625630630631u,0 563.063563063063u,1.5 564.0401031031031u,1.5 564.0411031031031u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 569.9053433433434u,0 569.9063433433433u,1.5 602.1641646646647u,1.5 602.1651646646646u,0 603.1417047047047u,0 603.1427047047047u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 606.0743248248249u,0 606.0753248248249u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 637.355606106106u,0 637.356606106106u,1.5 660.816567067067u,1.5 660.817567067067u,0 661.7941071071072u,0 661.7951071071071u,1.5 662.7716471471472u,1.5 662.7726471471472u,0 663.7491871871872u,0 663.7501871871872u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 685.255068068068u,0 685.256068068068u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 707.7384889889889u,1.5 707.7394889889889u,0 708.716029029029u,0 708.7170290290289u,1.5 709.693569069069u,1.5 709.694569069069u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 729.24436986987u,0 729.2453698698699u,1.5 730.22190990991u,1.5 730.22290990991u,0 731.19944994995u,0 731.20044994995u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 770.3010515515515u,0 770.3020515515515u,1.5 771.2785915915915u,1.5 771.2795915915915u,0 772.2561316316315u,0 772.2571316316315u,1.5 790.8293923923924u,1.5 790.8303923923924u,0 792.7844724724725u,0 792.7854724724725u,1.5 793.7620125125126u,1.5 793.7630125125125u,0 814.2903533533533u,0 814.2913533533533u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 816.2454334334335u,0 816.2464334334335u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 841.6614744744745u,1.5 841.6624744744745u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 868.0550555555556u,1.5 868.0560555555555u,0 869.0325955955957u,0 869.0335955955957u,1.5 894.4486366366367u,1.5 894.4496366366367u,0 896.4037167167166u,0 896.4047167167166u,1.5 897.3812567567567u,1.5 897.3822567567566u,0 927.684997997998u,0 927.685997997998u,1.5 928.6625380380381u,1.5 928.663538038038u,0 932.5726981981983u,0 932.5736981981983u,1.5 933.5502382382382u,1.5 933.5512382382382u,0 935.5053183183182u,0 935.5063183183182u,1.5 938.4379384384384u,1.5 938.4389384384384u,0 939.4154784784785u,0 939.4164784784784u,1.5 1057.6978233233233u,1.5 1057.6988233233235u,0 1058.6753633633632u,0 1058.6763633633634u,1.5 1061.6079834834834u,1.5 1061.6089834834836u,0 1062.5855235235235u,0 1062.5865235235237u,1.5 1065.5181436436435u,1.5 1065.5191436436437u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1070.4058438438437u,0 1070.406843843844u,1.5 1071.3833838838837u,1.5 1071.3843838838839u,0 1102.6646651651652u,0 1102.6656651651654u,1.5 1103.642205205205u,1.5 1103.6432052052053u,0 1104.6197452452452u,0 1104.6207452452454u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1107.5523653653654u,0 1107.5533653653656u,1.5 1108.5299054054053u,1.5 1108.5309054054055u,0 1109.5074454454455u,0 1109.5084454454457u,1.5 1134.9234864864864u,1.5 1134.9244864864866u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1161.3170675675676u,0 1161.3180675675678u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1163.2721476476477u,0 1163.2731476476479u,1.5 1164.2496876876876u,1.5 1164.2506876876878u,0 1165.2272277277275u,0 1165.2282277277277u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1208.2389894894895u,1.5 1208.2399894894897u,0 1210.1940695695696u,0 1210.1950695695698u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1231.6999504504504u,1.5 1231.7009504504506u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1254.1833713713713u,0 1254.1843713713715u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1269.8240120120117u,0 1269.825012012012u,1.5 1270.8015520520519u,1.5 1270.802552052052u,0 1271.779092092092u,0 1271.7800920920922u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1291.3298928928928u,1.5 1291.330892892893u,0 1292.3074329329327u,0 1292.3084329329329u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1315.7683938938937u,0 1315.769393893894u,1.5 1316.7459339339337u,1.5 1316.7469339339339u,0 1338.251814814815u,0 1338.252814814815u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1342.1619749749748u,0 1342.162974974975u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1367.578016016016u,0 1367.579016016016u,1.5 1368.5555560560558u,1.5 1368.556556056056u,0 1392.016517017017u,0 1392.017517017017u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1400.8143773773772u,1.5 1400.8153773773774u,0 1401.7919174174174u,0 1401.7929174174176u,1.5 1431.1181186186186u,1.5 1431.1191186186188u,0 1432.0956586586585u,0 1432.0966586586587u,1.5 1433.0731986986987u,1.5 1433.0741986986989u,0 1434.0507387387386u,0 1434.0517387387388u,1.5 1436.0058188188189u,1.5 1436.006818818819u,0 1438.938438938939u,0 1438.9394389389392u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1562.108483983984u,0 1562.109483983984u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1565.041104104104u,0 1565.0421041041043u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1567.973724224224u,0 1567.9747242242242u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1603.1651656656657u,0 1603.1661656656659u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1607.0753258258258u,1.5 1607.076325825826u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1662.795108108108u,1.5 1662.7961081081082u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1689.1886891891893u,1.5 1689.1896891891895u,0 1690.1662292292292u,0 1690.1672292292294u,1.5 1704.8293298298297u,1.5 1704.83032982983u,0 1705.8068698698698u,0 1705.80786986987u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1728.2902907907908u,0 1728.291290790791u,1.5 1729.2678308308307u,1.5 1729.268830830831u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1752.7287917917918u,1.5 1752.729791791792u,0 1767.3918923923923u,0 1767.3928923923925u,1.5 1768.3694324324322u,1.5 1768.3704324324324u,0 1771.3020525525524u,0 1771.3030525525526u,1.5 1790.852853353353u,1.5 1790.8538533533533u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1794.7630135135132u,0 1794.7640135135134u,1.5 1795.7405535535534u,1.5 1795.7415535535536u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1839.7298553553553u,1.5 1839.7308553553555u,0 1863.1908163163164u,0 1863.1918163163166u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1866.1234364364361u,0 1866.1244364364363u,1.5 1889.5843973973974u,1.5 1889.5853973973976u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1896.4271776776775u,1.5 1896.4281776776777u,0 1897.4047177177176u,0 1897.4057177177178u,1.5 1898.3822577577575u,1.5 1898.3832577577577u,0 1899.3597977977977u,0 1899.3607977977979u,1.5 1900.3373378378376u,1.5 1900.3383378378378u,0 1929.6635390390388u,0 1929.664539039039u,1.5 1930.641079079079u,1.5 1930.6420790790792u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1940.4164794794794u,1.5 1940.4174794794797u,0 1941.3940195195194u,0 1941.3950195195196u,1.5 1943.3490995995994u,1.5 1943.3500995995996u,0 1944.3266396396396u,0 1944.3276396396398u,1.5 2059.676364364364u,1.5 2059.677364364364u,0 2060.6539044044043u,0 2060.6549044044045u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2067.4966846846846u,1.5 2067.497684684685u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2070.429304804805u,1.5 2070.430304804805u,0 2103.665666166166u,0 2103.666666166166u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2105.620746246246u,0 2105.6217462462464u,1.5 2134.946947447447u,1.5 2134.9479474474474u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2137.8795675675674u,1.5 2137.8805675675676u,0 2138.8571076076073u,0 2138.8581076076075u,1.5 2139.8346476476477u,1.5 2139.835647647648u,0 2162.3180685685684u,0 2162.3190685685686u,1.5 2163.2956086086083u,1.5 2163.2966086086085u,0 2164.2731486486487u,0 2164.274148648649u,1.5 2184.8014894894895u,1.5 2184.8024894894897u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2187.7341096096093u,1.5 2187.7351096096095u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2227.813251251251u,1.5 2227.8142512512513u,0 2228.790791291291u,0 2228.7917912912912u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2230.745871371371u,0 2230.746871371371u,1.5 2231.7234114114112u,1.5 2231.7244114114114u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2254.2068323323324u,0 2254.2078323323326u,1.5 2268.869932932933u,1.5 2268.870932932933u,0 2269.847472972973u,0 2269.848472972973u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2290.3758138138137u,0 2290.376813813814u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2293.308433933934u,0 2293.309433933934u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2314.8143148148147u,0 2314.815314814815u,1.5 2316.769394894895u,1.5 2316.770394894895u,0 2317.746934934935u,0 2317.747934934935u,1.5 2318.724474974975u,1.5 2318.725474974975u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2340.2303558558556u,1.5 2340.231355855856u,0 2341.207895895896u,0 2341.208895895896u,1.5 2359.7811566566565u,1.5 2359.7821566566568u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2365.646396896897u,1.5 2365.647396896897u,0 2367.6014769769768u,0 2367.602476976977u,1.5 2368.5790170170167u,1.5 2368.580017017017u,0 2393.995058058058u,0 2393.996058058058u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2397.905218218218u,0 2397.9062182182183u,1.5 2432.119119619619u,1.5 2432.1201196196193u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2435.05173973974u,0 2435.05273973974u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.9843598598595u,0 2437.9853598598597u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2554.3116246246245u,0 2554.3126246246247u,1.5 2555.2891646646644u,1.5 2555.2901646646646u,0 2558.2217847847846u,0 2558.222784784785u,1.5 2559.1993248248245u,1.5 2559.2003248248247u,0 2560.1768648648645u,0 2560.1778648648647u,1.5 2562.1319449449447u,1.5 2562.132944944945u,0 2565.064565065065u,0 2565.065565065065u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2567.019645145145u,0 2567.0206451451454u,1.5 2567.997185185185u,1.5 2567.9981851851853u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2608.0763268268265u,1.5 2608.0773268268267u,0 2634.469907907908u,0 2634.470907907908u,1.5 2635.4474479479477u,1.5 2635.448447947948u,0 2637.402528028028u,0 2637.403528028028u,1.5 2657.9308688688684u,1.5 2657.9318688688686u,0 2658.9084089089088u,0 2658.909408908909u,1.5 2659.8859489489487u,1.5 2659.886948948949u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2665.751189189189u,0 2665.7521891891893u,1.5 2666.7287292292294u,1.5 2666.7297292292296u,0 2685.30198998999u,0 2685.3029899899902u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2689.21215015015u,1.5 2689.2131501501503u,0 2690.18969019019u,0 2690.1906901901903u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2710.718031031031u,0 2710.719031031031u,1.5 2711.695571071071u,1.5 2711.696571071071u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2730.268831831832u,0 2730.269831831832u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2750.7971726726723u,1.5 2750.7981726726725u,0 2751.7747127127127u,0 2751.775712712713u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2773.2805935935935u,0 2773.2815935935937u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2814.337275275275u,0 2814.338275275275u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2839.753316316316u,0 2839.7543163163164u,1.5 2840.730856356356u,1.5 2840.7318563563563u,0 2860.281657157157u,0 2860.2826571571572u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2865.169357357357u,1.5 2865.1703573573573u,0 2866.1468973973974u,0 2866.1478973973976u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2930.66454004004u,0 2930.66554004004u,1.5 2931.64208008008u,1.5 2931.6430800800804u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2938.48486036036u,1.5 2938.48586036036u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2941.4174804804807u,0 2941.418480480481u,1.5 2942.39502052052u,1.5 2942.3960205205203u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 3062.6324454454452u,1.5 3062.6334454454454u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3066.5426056056053u,0 3066.5436056056055u,1.5 3067.5201456456457u,1.5 3067.521145645646u,0 3103.689127127127u,0 3103.690127127127u,1.5 3104.666667167167u,1.5 3104.667667167167u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3135.947948448448u,1.5 3135.9489484484484u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3207.308371371371u,0 3207.309371371371u,1.5 3227.836712212212u,1.5 3227.8377122122124u,0 3228.814252252252u,0 3228.8152522522523u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3232.724412412412u,0 3232.7254124124124u,1.5 3233.701952452452u,1.5 3233.7029524524523u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3273.781094094094u,1.5 3273.782094094094u,0 3290.3992747747743u,0 3290.4002747747745u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3294.309434934935u,0 3294.310434934935u,1.5 3309.9500755755753u,1.5 3309.9510755755755u,0 3310.927615615615u,0 3310.9286156156154u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3335.366116616616u,0 3335.3671166166164u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3365.6698578578576u,0 3365.6708578578578u,1.5 3366.647397897898u,1.5 3366.648397897898u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3390.1083588588585u,1.5 3390.1093588588587u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3396.9511391391393u,0 3396.9521391391395u,1.5 3431.1650405405403u,1.5 3431.1660405405405u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3434.0976606606605u,1.5 3434.0986606606607u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3436.052740740741u,1.5 3436.053740740741u,0 3562.155405905906u,0 3562.156405905906u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.020646146146u,1.5 3568.0216461461464u,0 3568.998186186186u,0 3568.9991861861863u,1.5 3603.2120875875876u,1.5 3603.213087587588u,0 3605.1671676676674u,0 3605.1681676676676u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3607.1222477477477u,0 3607.123247747748u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3635.4709089089088u,0 3635.471908908909u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3637.425988988989u,0 3637.4269889889893u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3688.258071071071u,0 3688.259071071071u,1.5 3706.831331831832u,1.5 3706.832331831832u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3730.292292792793u,0 3730.293292792793u,1.5 3732.2473728728723u,1.5 3732.2483728728726u,0 3733.2249129129127u,0 3733.225912912913u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3772.326514514514u,0 3772.3275145145144u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3812.405656156156u,0 3812.4066561561563u,1.5 3813.383196196196u,1.5 3813.384196196196u,0 3814.3607362362363u,0 3814.3617362362365u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3816.315816316316u,0 3816.3168163163164u,1.5 3817.293356356356u,1.5 3817.2943563563563u,0 3818.2708963963964u,0 3818.2718963963966u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3836.844157157157u,0 3836.8451571571572u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3887.6762392392393u,1.5 3887.6772392392395u,0 3888.653779279279u,0 3888.6547792792794u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3895.4965595595595u,1.5 3895.4975595595597u,0 3933.6206211211206u,0 3933.621621121121u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3938.508321321321u,1.5 3938.5093213213213u,0 3939.4858613613615u,0 3939.4868613613617u,1.5 4057.768206206206u,1.5 4057.769206206206u,0 4058.7457462462457u,0 4058.746746246246u,1.5 4061.6783663663664u,1.5 4061.6793663663666u,0 4062.6559064064063u,0 4062.6569064064065u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4065.588526526526u,0 4065.5895265265262u,1.5 4066.566066566567u,1.5 4066.567066566567u,0 4067.5436066066063u,0 4067.5446066066065u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4101.757508008008u,0 4101.758508008008u,1.5 4102.735048048047u,1.5 4102.736048048047u,0 4104.690128128128u,0 4104.691128128128u,1.5 4105.667668168168u,1.5 4105.668668168169u,0 4106.645208208208u,0 4106.646208208208u,1.5 4134.993869369369u,1.5 4134.99486936937u,0 4137.9264894894895u,0 4137.92748948949u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4161.38745045045u,0 4161.38845045045u,1.5 4183.870871371371u,1.5 4183.8718713713715u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4209.286912412412u,0 4209.287912412412u,1.5 4225.9050930930935u,1.5 4225.906093093094u,0 4226.882633133133u,0 4226.883633133133u,1.5 4229.815253253253u,1.5 4229.816253253253u,0 4251.321134134134u,0 4251.322134134134u,1.5 4268.916854854855u,1.5 4268.917854854855u,0 4270.871934934935u,0 4270.872934934935u,1.5 4272.827015015015u,1.5 4272.828015015015u,0 4289.4451956956955u,0 4289.446195695696u,1.5 4290.422735735735u,1.5 4290.423735735735u,0 4292.377815815816u,0 4292.378815815816u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4294.3328958958955u,0 4294.333895895896u,1.5 4313.8836966966965u,1.5 4313.884696696697u,0 4336.367117617618u,0 4336.368117617618u,1.5 4337.344657657658u,1.5 4337.345657657658u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4342.232357857858u,0 4342.233357857858u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4362.760698698698u,0 4362.761698698699u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4368.625938938939u,0 4368.626938938939u,1.5 4369.603478978979u,1.5 4369.604478978979u,0 4390.13181981982u,0 4390.13281981982u,1.5 4391.10935985986u,1.5 4391.11035985986u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.99706006006u,0 4395.99806006006u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4438.031281781782u,1.5 4438.032281781782u,0 4440.963901901901u,0 4440.964901901902u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4565.111486986987u,0 4565.112486986987u,1.5 4566.0890270270265u,1.5 4566.090027027027u,0 4567.066567067067u,0 4567.067567067067u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4609.100788788789u,0 4609.101788788789u,1.5 4610.0783288288285u,1.5 4610.079328828829u,0 4635.49436986987u,0 4635.49536986987u,1.5 4636.471909909909u,1.5 4636.4729099099095u,0 4637.44944994995u,0 4637.45044994995u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4686.326451951952u,0 4686.327451951952u,1.5 4704.899712712712u,1.5 4704.900712712712u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4731.293293793794u,1.5 4731.294293793794u,0 4732.270833833833u,0 4732.271833833834u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4768.439815315315u,0 4768.440815315315u,1.5 4769.4173553553555u,1.5 4769.418355355356u,0 4771.372435435435u,0 4771.373435435436u,1.5 4793.8558563563565u,1.5 4793.856856356357u,0 4815.361737237236u,0 4815.362737237237u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4840.777778278279u,0 4840.778778278279u,1.5 4841.755318318318u,1.5 4841.756318318318u,0 4863.261199199199u,0 4863.262199199199u,1.5 4864.238739239238u,1.5 4864.239739239239u,0 4866.193819319319u,0 4866.194819319319u,1.5 4891.6098603603605u,1.5 4891.610860360361u,0 4892.5874004004u,0 4892.5884004004u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4894.542480480481u,0 4894.543480480481u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4898.45264064064u,0 4898.4536406406405u,1.5 4899.430180680681u,1.5 4899.431180680681u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4938.531782282283u,0 4938.532782282283u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 4941.464402402402u,0 4941.465402402402u,1.5 5057.791667167167u,1.5 5057.792667167168u,0 5058.769207207207u,0 5058.770207207207u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5064.634447447447u,1.5 5064.635447447447u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5135.99487037037u,0 5135.9958703703705u,1.5 5136.97241041041u,1.5 5136.97341041041u,0 5160.433371371371u,0 5160.4343713713715u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5162.388451451451u,0 5162.389451451451u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5208.332833333333u,0 5208.333833333333u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5232.771334334334u,1.5 5232.772334334334u,0 5250.367055055054u,0 5250.368055055054u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5289.468656656657u,0 5289.469656656657u,1.5 5290.4461966966965u,1.5 5290.447196696697u,0 5292.401276776777u,0 5292.402276776777u,1.5 5294.356356856857u,1.5 5294.357356856857u,0 5295.3338968968965u,0 5295.334896896897u,1.5 5312.929617617618u,1.5 5312.930617617618u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5337.368118618619u,0 5337.369118618619u,1.5 5338.345658658659u,1.5 5338.346658658659u,0 5339.323198698698u,0 5339.324198698699u,1.5 5362.78415965966u,1.5 5362.78515965966u,0 5363.761699699699u,0 5363.7626996997u,1.5 5364.739239739739u,1.5 5364.740239739739u,0 5366.69431981982u,0 5366.69531981982u,1.5 5367.67185985986u,1.5 5367.67285985986u,0 5394.065440940941u,0 5394.066440940941u,1.5 5395.042980980981u,1.5 5395.043980980981u,0 5396.020521021021u,0 5396.021521021021u,1.5 5396.998061061061u,1.5 5396.999061061061u,0 5397.975601101101u,0 5397.976601101102u,1.5 5398.953141141141u,1.5 5398.954141141141u,0 5399.930681181181u,0 5399.931681181181u,1.5 5430.2344224224225u,1.5 5430.235422422423u,0 5431.211962462463u,0 5431.212962462463u,1.5 5432.189502502502u,1.5 5432.190502502503u,0 5433.167042542542u,0 5433.168042542542u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5438.054742742742u,0 5438.055742742742u,1.5 5439.032282782783u,1.5 5439.033282782783u,0 5440.009822822823u,0 5440.010822822823u,1.5 5440.987362862863u,1.5 5440.988362862863u,0 5444.897523023023u,0 5444.898523023023u,1.5 5445.875063063063u,1.5 5445.876063063063u,0 5558.292167667668u,0 5558.293167667668u,1.5 5559.269707707707u,1.5 5559.2707077077075u,0 5562.2023278278275u,0 5562.203327827828u,1.5 5563.179867867868u,1.5 5563.180867867868u,0 5566.112487987988u,0 5566.113487987988u,1.5 5567.0900280280275u,1.5 5567.091028028028u,0 5568.067568068068u,0 5568.068568068068u,1.5 5570.022648148148u,1.5 5570.023648148148u,0 5571.000188188188u,0 5571.001188188188u,1.5 5600.326389389389u,1.5 5600.327389389389u,0 5601.303929429429u,0 5601.30492942943u,1.5 5605.21408958959u,1.5 5605.21508958959u,0 5608.146709709709u,0 5608.1477097097095u,1.5 5609.12424974975u,1.5 5609.12524974975u,0 5633.562750750751u,0 5633.563750750751u,1.5 5634.540290790791u,1.5 5634.541290790791u,0 5636.495370870871u,0 5636.496370870871u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5638.450450950951u,0 5638.451450950951u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5664.8440320320315u,0 5664.845032032032u,1.5 5665.821572072072u,1.5 5665.822572072072u,0 5682.439752752753u,0 5682.440752752753u,1.5 5683.417292792793u,1.5 5683.418292792793u,0 5685.372372872873u,0 5685.373372872873u,1.5 5688.304992992993u,1.5 5688.305992992993u,0 5689.282533033032u,0 5689.283533033033u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5727.406594594595u,0 5727.407594594595u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5772.373436436436u,0 5772.374436436437u,1.5 5788.991617117117u,1.5 5788.992617117117u,0 5789.9691571571575u,0 5789.970157157158u,1.5 5790.946697197197u,1.5 5790.947697197197u,0 5792.901777277278u,0 5792.902777277278u,1.5 5793.879317317317u,1.5 5793.880317317317u,0 5813.430118118118u,0 5813.431118118118u,1.5 5815.385198198198u,1.5 5815.386198198198u,0 5816.362738238237u,0 5816.363738238238u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5838.8461591591595u,0 5838.84715915916u,1.5 5840.801239239238u,1.5 5840.802239239239u,0 5859.3745u,0 5859.3755u,1.5 5860.352040040039u,1.5 5860.35304004004u,0 5862.30712012012u,0 5862.30812012012u,1.5 5863.2846601601605u,1.5 5863.285660160161u,0 5864.2622002002u,0 5864.2632002002u,1.5 5888.700701201201u,1.5 5888.701701201201u,0 5889.67824124124u,0 5889.679241241241u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5899.453641641641u,0 5899.4546416416415u,1.5 5900.431181681682u,1.5 5900.432181681682u,0 5932.690003003003u,0 5932.691003003003u,1.5 5933.667543043042u,1.5 5933.6685430430425u,0 5935.622623123123u,0 5935.623623123123u,1.5 5936.600163163163u,1.5 5936.601163163164u,0 5938.555243243242u,0 5938.5562432432425u,1.5 6055.860048048047u,1.5 6055.861048048047u,0 6056.8375880880885u,0 6056.838588088089u,1.5 6059.770208208208u,1.5 6059.771208208208u,0 6060.747748248248u,0 6060.748748248248u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6068.568068568568u,0 6068.569068568569u,1.5 6070.523148648648u,1.5 6070.524148648648u,0 6071.500688688689u,0 6071.501688688689u,1.5 6072.478228728728u,1.5 6072.479228728728u,0 6074.433308808809u,0 6074.434308808809u,1.5 6075.410848848848u,1.5 6075.411848848848u,0 6101.80442992993u,0 6101.80542992993u,1.5 6102.78196996997u,1.5 6102.7829699699705u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6106.69213013013u,0 6106.69313013013u,1.5 6107.66967017017u,1.5 6107.6706701701705u,0 6108.64721021021u,0 6108.64821021021u,1.5 6136.018331331331u,1.5 6136.019331331331u,0 6137.973411411411u,0 6137.974411411411u,1.5 6138.950951451451u,1.5 6138.951951451451u,0 6139.9284914914915u,0 6139.929491491492u,1.5 6140.906031531531u,1.5 6140.907031531531u,0 6159.4792922922925u,0 6159.480292292293u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6162.411912412412u,0 6162.412912412412u,1.5 6184.895333333333u,1.5 6184.896333333333u,0 6185.872873373373u,0 6185.8738733733735u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6208.3562942942945u,0 6208.357294294295u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6231.817255255255u,0 6231.818255255255u,1.5 6232.794795295295u,1.5 6232.795795295296u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6268.963776776777u,1.5 6268.964776776777u,0 6269.941316816817u,0 6269.942316816817u,1.5 6270.918856856857u,1.5 6270.919856856857u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6272.873936936937u,1.5 6272.874936936937u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6291.447197697697u,0 6291.448197697698u,1.5 6313.930618618619u,1.5 6313.931618618619u,0 6314.908158658659u,0 6314.909158658659u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6317.840778778779u,0 6317.841778778779u,1.5 6318.818318818819u,1.5 6318.819318818819u,0 6337.391579579579u,0 6337.392579579579u,1.5 6339.34665965966u,1.5 6339.34765965966u,0 6340.324199699699u,0 6340.3251996997u,1.5 6342.27927977978u,1.5 6342.28027977978u,0 6343.25681981982u,0 6343.25781981982u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6363.785160660661u,1.5 6363.786160660661u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6397.021522022022u,0 6397.022522022022u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6437.100663663664u,1.5 6437.101663663664u,0 6446.876064064064u,0 6446.877064064064u,1.5 6447.853604104104u,1.5 6447.8546041041045u,0 6562.225788788789u,0 6562.226788788789u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6565.158408908908u,1.5 6565.1594089089085u,0 6566.135948948949u,0 6566.136948948949u,1.5 6568.0910290290285u,1.5 6568.092029029029u,0 6569.068569069069u,0 6569.069569069069u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.001189189189u,0 6572.002189189189u,1.5 6600.34985035035u,1.5 6600.35085035035u,0 6601.32739039039u,0 6601.32839039039u,1.5 6604.26001051051u,1.5 6604.2610105105105u,0 6606.215090590591u,0 6606.216090590591u,1.5 6607.19263063063u,1.5 6607.193630630631u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6637.496371871872u,0 6637.497371871872u,1.5 6638.473911911911u,1.5 6638.4749119119115u,0 6639.451451951952u,0 6639.452451951952u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6664.867492992993u,0 6664.868492992993u,1.5 6665.845033033032u,1.5 6665.846033033033u,0 6685.395833833833u,0 6685.396833833834u,1.5 6705.924174674675u,1.5 6705.925174674675u,0 6706.901714714714u,0 6706.902714714714u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6708.856794794795u,0 6708.857794794795u,1.5 6709.834334834834u,1.5 6709.835334834835u,0 6726.452515515515u,0 6726.453515515515u,1.5 6727.430055555555u,1.5 6727.431055555555u,0 6729.385135635635u,0 6729.386135635636u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6752.846096596597u,1.5 6752.847096596597u,0 6768.486737237236u,0 6768.487737237237u,1.5 6769.464277277278u,1.5 6769.465277277278u,0 6771.4193573573575u,0 6771.420357357358u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6791.947698198198u,1.5 6791.948698198198u,0 6813.453579079079u,0 6813.454579079079u,1.5 6814.431119119119u,1.5 6814.432119119119u,0 6815.4086591591595u,0 6815.40965915916u,1.5 6835.937u,1.5 6835.938u,0 6837.89208008008u,0 6837.89308008008u,1.5 6839.8471601601605u,1.5 6839.848160160161u,0 6860.375501001001u,0 6860.376501001001u,1.5 6861.35304104104u,1.5 6861.354041041041u,0 6864.285661161161u,0 6864.286661161162u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6867.218281281282u,0 6867.219281281282u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6893.611862362362u,0 6893.612862362363u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6932.713463963964u,0 6932.714463963965u,1.5 6933.691004004004u,1.5 6933.692004004004u,0 6934.668544044043u,0 6934.6695440440435u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6936.623624124124u,0 6936.624624124124u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6939.556244244243u,0 6939.5572442442435u,1.5 6942.488864364364u,1.5 6942.489864364365u,0 6943.466404404404u,0 6943.467404404404u,1.5
vbb14 bb14 0 pwl 0,1.5  104.59628428428428u,1.5 104.59728428428429u,0 106.55136436436436u,0 106.55236436436437u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 109.48398448448448u,0 109.48498448448449u,1.5 110.46152452452452u,1.5 110.46252452452453u,0 158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 164.22622672672674u,0 164.2272267267267u,1.5 207.2379884884885u,1.5 207.23898848848847u,0 208.21552852852852u,0 208.2165285285285u,1.5 210.17060860860863u,1.5 210.1716086086086u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 289.35135185185186u,1.5 289.35235185185184u,0 290.32889189189194u,0 290.3298918918919u,1.5 294.23905205205205u,1.5 294.240052052052u,0 335.2957337337337u,0 335.2967337337337u,1.5 336.2732737737738u,1.5 336.27427377377376u,0 337.2508138138138u,0 337.2518138138138u,1.5 338.2283538538539u,1.5 338.22935385385387u,0 340.18343393393394u,0 340.1844339339339u,1.5 389.06043593593597u,1.5 389.06143593593595u,0 390.037975975976u,0 390.038975975976u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 395.90321621621626u,1.5 395.90421621621624u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 602.1641646646647u,0 602.1651646646646u,1.5 603.1417047047047u,1.5 603.1427047047047u,0 605.0967847847849u,0 605.0977847847848u,1.5 606.0743248248249u,1.5 606.0753248248249u,0 607.0518648648649u,0 607.0528648648649u,1.5 660.816567067067u,1.5 660.817567067067u,0 661.7941071071072u,0 661.7951071071071u,1.5 662.7716471471472u,1.5 662.7726471471472u,0 663.7491871871872u,0 663.7501871871872u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 707.7384889889889u,0 707.7394889889889u,1.5 708.716029029029u,1.5 708.7170290290289u,0 709.693569069069u,0 709.694569069069u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 790.8293923923924u,0 790.8303923923924u,1.5 792.7844724724725u,1.5 792.7854724724725u,0 793.7620125125126u,0 793.7630125125125u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 841.6614744744745u,1.5 841.6624744744745u,0 894.4486366366367u,0 894.4496366366367u,1.5 896.4037167167166u,1.5 896.4047167167166u,0 897.3812567567567u,0 897.3822567567566u,1.5 1102.6646651651652u,1.5 1102.6656651651654u,0 1103.642205205205u,0 1103.6432052052053u,1.5 1104.6197452452452u,1.5 1104.6207452452454u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1107.5523653653654u,1.5 1107.5533653653656u,0 1108.5299054054053u,0 1108.5309054054055u,1.5 1109.5074454454455u,1.5 1109.5084454454457u,0 1161.3170675675676u,0 1161.3180675675678u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1163.2721476476477u,0 1163.2731476476479u,1.5 1164.2496876876876u,1.5 1164.2506876876878u,0 1165.2272277277275u,0 1165.2282277277277u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1208.2389894894895u,0 1208.2399894894897u,1.5 1210.1940695695696u,1.5 1210.1950695695698u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1254.1833713713713u,0 1254.1843713713715u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1291.3298928928928u,0 1291.330892892893u,1.5 1292.3074329329327u,1.5 1292.3084329329329u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1338.251814814815u,0 1338.252814814815u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1342.1619749749748u,0 1342.162974974975u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1400.8143773773772u,0 1400.8153773773774u,1.5 1401.7919174174174u,1.5 1401.7929174174176u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1603.1651656656657u,1.5 1603.1661656656659u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1607.0753258258258u,0 1607.076325825826u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1662.795108108108u,1.5 1662.7961081081082u,0 1704.8293298298297u,0 1704.83032982983u,1.5 1705.8068698698698u,1.5 1705.80786986987u,0 1707.76194994995u,0 1707.76294994995u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1752.7287917917918u,1.5 1752.729791791792u,0 1790.852853353353u,0 1790.8538533533533u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1794.7630135135132u,1.5 1794.7640135135134u,0 1795.7405535535534u,0 1795.7415535535536u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1839.7298553553553u,1.5 1839.7308553553555u,0 1889.5843973973974u,0 1889.5853973973976u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1896.4271776776775u,0 1896.4281776776777u,1.5 1897.4047177177176u,1.5 1897.4057177177178u,0 1898.3822577577575u,0 1898.3832577577577u,1.5 1899.3597977977977u,1.5 1899.3607977977979u,0 1900.3373378378376u,0 1900.3383378378378u,1.5 2103.665666166166u,1.5 2103.666666166166u,0 2104.643206206206u,0 2104.644206206206u,1.5 2105.620746246246u,1.5 2105.6217462462464u,0 2162.3180685685684u,0 2162.3190685685686u,1.5 2163.2956086086083u,1.5 2163.2966086086085u,0 2164.2731486486487u,0 2164.274148648649u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2254.2068323323324u,0 2254.2078323323326u,1.5 2290.3758138138137u,1.5 2290.376813813814u,0 2292.330893893894u,0 2292.331893893894u,1.5 2293.308433933934u,1.5 2293.309433933934u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2340.2303558558556u,1.5 2340.231355855856u,0 2341.207895895896u,0 2341.208895895896u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2397.905218218218u,1.5 2397.9062182182183u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2608.0763268268265u,0 2608.0773268268267u,1.5 2657.9308688688684u,1.5 2657.9318688688686u,0 2658.9084089089088u,0 2658.909408908909u,1.5 2659.8859489489487u,1.5 2659.886948948949u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2665.751189189189u,0 2665.7521891891893u,1.5 2666.7287292292294u,1.5 2666.7297292292296u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2710.718031031031u,1.5 2710.719031031031u,0 2711.695571071071u,0 2711.696571071071u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2750.7971726726723u,1.5 2750.7981726726725u,0 2751.7747127127127u,0 2751.775712712713u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2839.753316316316u,0 2839.7543163163164u,1.5 2840.730856356356u,1.5 2840.7318563563563u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3104.666667167167u,0 3104.667667167167u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3207.308371371371u,1.5 3207.309371371371u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3290.3992747747743u,1.5 3290.4002747747745u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3294.309434934935u,1.5 3294.310434934935u,0 3335.366116616616u,0 3335.3671166166164u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3390.1083588588585u,0 3390.1093588588587u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.996059059059u,0 3394.997059059059u,1.5 3396.9511391391393u,1.5 3396.9521391391395u,0 3603.2120875875876u,0 3603.213087587588u,1.5 3605.1671676676674u,1.5 3605.1681676676676u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3607.1222477477477u,1.5 3607.123247747748u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3706.831331831832u,0 3706.832331831832u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3836.844157157157u,0 3836.8451571571572u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 3887.6762392392393u,0 3887.6772392392395u,1.5 3888.653779279279u,1.5 3888.6547792792794u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3895.4965595595595u,0 3895.4975595595597u,1.5 4101.757508008008u,1.5 4101.758508008008u,0 4102.735048048047u,0 4102.736048048047u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4105.667668168168u,0 4105.668668168169u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4161.38745045045u,0 4161.38845045045u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4209.286912412412u,1.5 4209.287912412412u,0 4251.321134134134u,0 4251.322134134134u,1.5 4289.4451956956955u,1.5 4289.446195695696u,0 4290.422735735735u,0 4290.423735735735u,1.5 4292.377815815816u,1.5 4292.378815815816u,0 4293.355355855856u,0 4293.356355855856u,1.5 4294.3328958958955u,1.5 4294.333895895896u,0 4336.367117617618u,0 4336.368117617618u,1.5 4337.344657657658u,1.5 4337.345657657658u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4342.232357857858u,0 4342.233357857858u,1.5 4390.13181981982u,1.5 4390.13281981982u,0 4391.10935985986u,0 4391.11035985986u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.99706006006u,1.5 4395.99806006006u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4609.100788788789u,1.5 4609.101788788789u,0 4610.0783288288285u,0 4610.079328828829u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4704.899712712712u,0 4704.900712712712u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4793.8558563563565u,0 4793.856856356357u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4840.777778278279u,0 4840.778778278279u,1.5 4841.755318318318u,1.5 4841.756318318318u,0 4891.6098603603605u,0 4891.610860360361u,1.5 4892.5874004004u,1.5 4892.5884004004u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4894.542480480481u,1.5 4894.543480480481u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4898.45264064064u,1.5 4898.4536406406405u,0 4899.430180680681u,0 4899.431180680681u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5160.433371371371u,0 5160.4343713713715u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5162.388451451451u,0 5162.389451451451u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5250.367055055054u,0 5250.368055055054u,1.5 5289.468656656657u,1.5 5289.469656656657u,0 5290.4461966966965u,0 5290.447196696697u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5294.356356856857u,0 5294.357356856857u,1.5 5295.3338968968965u,1.5 5295.334896896897u,0 5337.368118618619u,0 5337.369118618619u,1.5 5338.345658658659u,1.5 5338.346658658659u,0 5339.323198698698u,0 5339.324198698699u,1.5 5394.065440940941u,1.5 5394.066440940941u,0 5395.042980980981u,0 5395.043980980981u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5396.998061061061u,0 5396.999061061061u,1.5 5397.975601101101u,1.5 5397.976601101102u,0 5398.953141141141u,0 5398.954141141141u,1.5 5399.930681181181u,1.5 5399.931681181181u,0 5600.326389389389u,0 5600.327389389389u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5605.21408958959u,0 5605.21508958959u,1.5 5608.146709709709u,1.5 5608.1477097097095u,0 5609.12424974975u,0 5609.12524974975u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5664.8440320320315u,0 5664.845032032032u,1.5 5665.821572072072u,1.5 5665.822572072072u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 5788.991617117117u,0 5788.992617117117u,1.5 5789.9691571571575u,1.5 5789.970157157158u,0 5790.946697197197u,0 5790.947697197197u,1.5 5792.901777277278u,1.5 5792.902777277278u,0 5793.879317317317u,0 5793.880317317317u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5838.8461591591595u,0 5838.84715915916u,1.5 5840.801239239238u,1.5 5840.802239239239u,0 5888.700701201201u,0 5888.701701201201u,1.5 5889.67824124124u,1.5 5889.679241241241u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5899.453641641641u,1.5 5899.4546416416415u,0 5900.431181681682u,0 5900.432181681682u,1.5 6101.80442992993u,1.5 6101.80542992993u,0 6102.78196996997u,0 6102.7829699699705u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6106.69213013013u,1.5 6106.69313013013u,0 6107.66967017017u,0 6107.6706701701705u,1.5 6108.64721021021u,1.5 6108.64821021021u,0 6159.4792922922925u,0 6159.480292292293u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6162.411912412412u,0 6162.412912412412u,1.5 6208.3562942942945u,1.5 6208.357294294295u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6291.447197697697u,1.5 6291.448197697698u,0 6337.391579579579u,0 6337.392579579579u,1.5 6339.34665965966u,1.5 6339.34765965966u,0 6340.324199699699u,0 6340.3251996997u,1.5 6342.27927977978u,1.5 6342.28027977978u,0 6343.25681981982u,0 6343.25781981982u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6600.34985035035u,0 6600.35085035035u,1.5 6601.32739039039u,1.5 6601.32839039039u,0 6604.26001051051u,0 6604.2610105105105u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6607.19263063063u,0 6607.193630630631u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6664.867492992993u,0 6664.868492992993u,1.5 6665.845033033032u,1.5 6665.846033033033u,0 6705.924174674675u,0 6705.925174674675u,1.5 6706.901714714714u,1.5 6706.902714714714u,0 6707.879254754755u,0 6707.880254754755u,1.5 6708.856794794795u,1.5 6708.857794794795u,0 6709.834334834834u,0 6709.835334834835u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6752.846096596597u,1.5 6752.847096596597u,0 6791.947698198198u,0 6791.948698198198u,1.5 6835.937u,1.5 6835.938u,0 6837.89208008008u,0 6837.89308008008u,1.5 6839.8471601601605u,1.5 6839.848160160161u,0 6892.634322322322u,0 6892.635322322322u,1.5 6893.611862362362u,1.5 6893.612862362363u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5
vbb15 bb15 0 pwl 0,1.5  158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 164.22622672672674u,1.5 164.2272267267267u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 336.2732737737738u,0 336.27427377377376u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 338.2283538538539u,0 338.22935385385387u,1.5 340.18343393393394u,1.5 340.1844339339339u,0 660.816567067067u,0 660.817567067067u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 662.7716471471472u,0 662.7726471471472u,1.5 663.7491871871872u,1.5 663.7501871871872u,0 664.7267272272272u,0 664.7277272272272u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 841.6614744744745u,0 841.6624744744745u,1.5 1161.3170675675676u,1.5 1161.3180675675678u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1163.2721476476477u,1.5 1163.2731476476479u,0 1164.2496876876876u,0 1164.2506876876878u,1.5 1165.2272277277275u,1.5 1165.2282277277277u,0 1249.295671171171u,0 1249.2966711711713u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1251.2507512512511u,0 1251.2517512512513u,1.5 1253.2058313313312u,1.5 1253.2068313313314u,0 1254.1833713713713u,0 1254.1843713713715u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1342.1619749749748u,1.5 1342.162974974975u,0 1662.795108108108u,0 1662.7961081081082u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1752.7287917917918u,1.5 1752.729791791792u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1839.7298553553553u,0 1839.7308553553555u,1.5 2162.3180685685684u,1.5 2162.3190685685686u,0 2163.2956086086083u,0 2163.2966086086085u,1.5 2164.2731486486487u,1.5 2164.274148648649u,0 2250.296672172172u,0 2250.297672172172u,1.5 2253.2292922922925u,1.5 2253.2302922922927u,0 2254.2068323323324u,0 2254.2078323323326u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2340.2303558558556u,0 2340.231355855856u,1.5 2341.207895895896u,1.5 2341.208895895896u,0 2657.9308688688684u,0 2657.9318688688686u,1.5 2658.9084089089088u,1.5 2658.909408908909u,0 2659.8859489489487u,0 2659.886948948949u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2665.751189189189u,1.5 2665.7521891891893u,0 2666.7287292292294u,0 2666.7297292292296u,1.5 2748.8420925925925u,1.5 2748.8430925925927u,0 2749.819632632633u,0 2749.820632632633u,1.5 2750.7971726726723u,1.5 2750.7981726726725u,0 2751.7747127127127u,0 2751.775712712713u,1.5 2752.7522527527526u,1.5 2752.753252752753u,0 2753.729792792793u,0 2753.730792792793u,1.5 2754.707332832833u,1.5 2754.708332832833u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2839.753316316316u,1.5 2839.7543163163164u,0 2840.730856356356u,0 2840.7318563563563u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3250.3201331331334u,0 3250.3211331331336u,1.5 3335.366116616616u,1.5 3335.3671166166164u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3836.844157157157u,1.5 3836.8451571571572u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4251.321134134134u,0 4251.322134134134u,1.5 4336.367117617618u,1.5 4336.368117617618u,0 4337.344657657658u,0 4337.345657657658u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4342.232357857858u,1.5 4342.233357857858u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4750.844094594595u,1.5 4750.845094594595u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4840.777778278279u,1.5 4840.778778278279u,0 4841.755318318318u,0 4841.756318318318u,1.5 5160.433371371371u,1.5 5160.4343713713715u,0 5161.410911411411u,0 5161.411911411411u,1.5 5162.388451451451u,1.5 5162.389451451451u,0 5250.367055055054u,0 5250.368055055054u,1.5 5337.368118618619u,1.5 5337.369118618619u,0 5338.345658658659u,0 5338.346658658659u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5664.8440320320315u,1.5 5664.845032032032u,0 5665.821572072072u,0 5665.822572072072u,1.5 5749.890015515515u,1.5 5749.891015515515u,0 5750.867555555555u,0 5750.868555555555u,1.5 5751.845095595596u,1.5 5751.846095595596u,0 5837.868619119119u,0 5837.869619119119u,1.5 5838.8461591591595u,1.5 5838.84715915916u,0 5840.801239239238u,0 5840.802239239239u,1.5 6159.4792922922925u,1.5 6159.480292292293u,0 6160.456832332332u,0 6160.457832332332u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6337.391579579579u,1.5 6337.392579579579u,0 6339.34665965966u,0 6339.34765965966u,1.5 6340.324199699699u,1.5 6340.3251996997u,0 6342.27927977978u,0 6342.28027977978u,1.5 6343.25681981982u,1.5 6343.25781981982u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6664.867492992993u,1.5 6664.868492992993u,0 6665.845033033032u,0 6665.846033033033u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6749.913476476477u,0 6749.914476476477u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6751.868556556556u,0 6751.869556556556u,1.5 6752.846096596597u,1.5 6752.847096596597u,0 6835.937u,0 6835.938u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6839.8471601601605u,0 6839.848160160161u,1.5
vbb16 bb16 0 pwl 0,1.5  249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 1249.295671171171u,1.5 1249.2966711711713u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1251.2507512512511u,1.5 1251.2517512512513u,0 1253.2058313313312u,0 1253.2068313313314u,1.5 1254.1833713713713u,1.5 1254.1843713713715u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1752.7287917917918u,0 1752.729791791792u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2253.2292922922925u,0 2253.2302922922927u,1.5 2254.2068323323324u,1.5 2254.2078323323326u,0 2748.8420925925925u,0 2748.8430925925927u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2750.7971726726723u,0 2750.7981726726725u,1.5 2751.7747127127127u,1.5 2751.775712712713u,0 2752.7522527527526u,0 2752.753252752753u,1.5 2753.729792792793u,1.5 2753.730792792793u,0 2754.707332832833u,0 2754.708332832833u,1.5 3250.3201331331334u,1.5 3250.3211331331336u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4750.844094594595u,0 4750.845094594595u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5749.890015515515u,0 5749.891015515515u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5751.845095595596u,0 5751.846095595596u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6748.935936436436u,0 6748.936936436437u,1.5 6749.913476476477u,1.5 6749.914476476477u,0 6750.891016516516u,0 6750.892016516516u,1.5 6751.868556556556u,1.5 6751.869556556556u,0 6752.846096596597u,0 6752.847096596597u,1.5

vb21 b21 0 pwl 0,1.5  2.93212012012012u,1.5 2.9331201201201202u,0 3.90966016016016u,0 3.9106601601601603u,1.5 10.75244044044044u,1.5 10.753440440440441u,0 11.72998048048048u,0 11.730980480480481u,1.5 17.59522072072072u,1.5 17.59622072072072u,0 18.572760760760765u,0 18.573760760760763u,1.5 21.50538088088088u,1.5 21.50638088088088u,0 22.482920920920925u,0 22.483920920920923u,1.5 27.370621121121122u,1.5 27.37162112112112u,0 28.348161161161162u,0 28.34916116116116u,1.5 29.325701201201202u,1.5 29.3267012012012u,0 30.303241241241246u,0 30.304241241241243u,1.5 32.25832132132132u,1.5 32.25932132132132u,0 37.146021521521526u,0 37.14702152152153u,1.5 38.12356156156156u,1.5 38.12456156156156u,0 40.07864164164164u,0 40.07964164164164u,1.5 41.05618168168168u,1.5 41.05718168168168u,0 42.03372172172172u,0 42.03472172172172u,1.5 43.01126176176176u,1.5 43.01226176176176u,0 46.92142192192192u,0 46.922421921921924u,1.5 47.89896196196196u,1.5 47.899961961961964u,0 49.85404204204204u,0 49.855042042042044u,1.5 51.80912212212212u,1.5 51.810122122122124u,0 52.786662162162166u,0 52.78766216216217u,1.5 56.69682232232232u,1.5 56.697822322322324u,0 57.67436236236236u,0 57.675362362362364u,1.5 61.58452252252251u,1.5 61.58552252252252u,0 62.56206256256256u,0 62.563062562562564u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 64.51714264264264u,0 64.51814264264264u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 67.44976276276276u,1.5 67.45076276276276u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 70.38238288288288u,0 70.38338288288288u,1.5 71.35992292292292u,1.5 71.36092292292292u,0 73.315003003003u,0 73.316003003003u,1.5 75.27008308308308u,1.5 75.27108308308308u,0 77.22516316316316u,0 77.22616316316316u,1.5 78.2027032032032u,1.5 78.2037032032032u,0 79.18024324324324u,0 79.18124324324324u,1.5 81.13532332332332u,1.5 81.13632332332332u,0 83.0904034034034u,0 83.0914034034034u,1.5 85.04548348348348u,1.5 85.04648348348348u,0 86.02302352352352u,0 86.02402352352352u,1.5 88.95564364364364u,1.5 88.95664364364364u,0 89.9331836836837u,0 89.9341836836837u,1.5 90.91072372372372u,1.5 90.91172372372372u,0 92.8658038038038u,0 92.8668038038038u,1.5 93.84334384384384u,1.5 93.84434384384384u,0 96.77596396396396u,0 96.77696396396396u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 114.37168468468468u,0 114.37268468468469u,1.5 115.34922472472472u,1.5 115.35022472472473u,0 116.32676476476476u,0 116.32776476476477u,1.5 120.23692492492492u,1.5 120.23792492492493u,0 121.21446496496498u,0 121.21546496496498u,1.5 122.19200500500502u,1.5 122.19300500500502u,0 124.14708508508508u,0 124.14808508508509u,1.5 125.12462512512512u,1.5 125.12562512512513u,0 129.0347852852853u,0 129.03578528528527u,1.5 130.01232532532532u,1.5 130.0133253253253u,0 130.98986536536538u,0 130.99086536536535u,1.5 134.90002552552554u,1.5 134.9010255255255u,0 135.8775655655656u,0 135.87856556556557u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 141.74280580580583u,0 141.7438058058058u,1.5 143.69788588588588u,1.5 143.69888588588586u,0 144.67542592592594u,0 144.6764259259259u,1.5 148.58558608608612u,1.5 148.5865860860861u,0 149.56312612612612u,0 149.5641261261261u,1.5 150.54066616616618u,1.5 150.54166616616615u,0 151.51820620620623u,0 151.5192062062062u,1.5 152.49574624624626u,1.5 152.49674624624623u,0 156.40590640640642u,0 156.4069064064064u,1.5 158.3609864864865u,1.5 158.36198648648647u,0 159.33852652652652u,0 159.3395265265265u,1.5 163.2486866866867u,1.5 163.2496866866867u,0 165.20376676676676u,0 165.20476676676674u,1.5 166.18130680680682u,1.5 166.1823068068068u,0 169.11392692692695u,0 169.11492692692693u,1.5 174.00162712712714u,1.5 174.0026271271271u,0 177.9117872872873u,0 177.91278728728727u,1.5 179.8668673673674u,1.5 179.86786736736738u,0 180.8444074074074u,0 180.84540740740738u,1.5 182.7994874874875u,1.5 182.8004874874875u,0 183.77702752752754u,0 183.7780275275275u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 190.6198078078078u,0 190.62080780780778u,1.5 192.57488788788788u,1.5 192.57588788788786u,0 193.55242792792794u,0 193.5534279279279u,1.5 194.529967967968u,1.5 194.53096796796797u,0 195.50750800800802u,0 195.508508008008u,1.5 197.4625880880881u,1.5 197.46358808808807u,0 201.37274824824826u,0 201.37374824824823u,1.5 203.32782832832834u,1.5 203.3288283283283u,0 204.3053683683684u,0 204.30636836836837u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 215.05830880880882u,0 215.0593088088088u,1.5 217.0133888888889u,1.5 217.01438888888887u,0 217.99092892892892u,0 217.9919289289289u,1.5 218.96846896896898u,1.5 218.96946896896895u,0 221.90108908908908u,0 221.90208908908906u,1.5 223.85616916916916u,1.5 223.85716916916914u,0 224.83370920920922u,0 224.8347092092092u,1.5 225.81124924924927u,1.5 225.81224924924925u,0 226.7887892892893u,0 226.78978928928927u,1.5 228.74386936936938u,1.5 228.74486936936935u,0 234.60910960960962u,0 234.6101096096096u,1.5 239.4968098098098u,1.5 239.49780980980978u,0 242.42942992992997u,0 242.43042992992994u,1.5 243.40696996996996u,1.5 243.40796996996994u,0 245.36205005005007u,0 245.36305005005005u,1.5 247.31713013013015u,1.5 247.31813013013013u,0 248.29467017017018u,0 248.29567017017015u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 255.13745045045044u,0 255.13845045045042u,1.5 259.04761061061066u,1.5 259.04861061061064u,0 260.02515065065063u,0 260.0261506506506u,1.5 261.98023073073074u,1.5 261.9812307307307u,0 262.95777077077076u,0 262.95877077077074u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 274.68825125125124u,0 274.6892512512512u,1.5 280.5534914914915u,1.5 280.5544914914915u,0 281.53103153153154u,0 281.5320315315315u,1.5 282.50857157157157u,1.5 282.50957157157154u,0 283.48611161161165u,0 283.4871116116116u,1.5 285.4411916916917u,1.5 285.4421916916917u,0 287.39627177177175u,0 287.3972717717717u,1.5 291.3064319319319u,1.5 291.3074319319319u,0 292.28397197197194u,0 292.2849719719719u,1.5 294.23905205205205u,1.5 294.240052052052u,0 299.12675225225223u,0 299.1277522522522u,1.5 302.0593723723724u,1.5 302.0603723723724u,0 303.03691241241245u,0 303.0379124124124u,1.5 304.9919924924925u,1.5 304.9929924924925u,0 305.9695325325325u,0 305.9705325325325u,1.5 306.9470725725726u,1.5 306.9480725725726u,0 308.90215265265266u,0 308.90315265265264u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 316.722472972973u,0 316.72347297297296u,1.5 317.700013013013u,1.5 317.701013013013u,0 318.67755305305303u,0 318.678553053053u,1.5 319.6550930930931u,1.5 319.6560930930931u,0 320.63263313313314u,0 320.6336331331331u,1.5 325.5203333333333u,1.5 325.5213333333333u,0 326.4978733733734u,0 326.4988733733734u,1.5 327.47541341341343u,1.5 327.4764134134134u,0 329.4304934934935u,0 329.43149349349346u,1.5 331.3855735735736u,1.5 331.38657357357357u,0 332.3631136136136u,0 332.3641136136136u,1.5 333.3406536536537u,1.5 333.3416536536537u,0 335.2957337337337u,0 335.2967337337337u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 342.138514014014u,0 342.13951401401397u,1.5 343.1160540540541u,1.5 343.11705405405405u,0 345.0711341341341u,0 345.0721341341341u,1.5 346.0486741741742u,1.5 346.0496741741742u,0 347.02621421421424u,0 347.0272142142142u,1.5 348.9812942942943u,1.5 348.98229429429426u,0 349.9588343343343u,0 349.9598343343343u,1.5 350.9363743743744u,1.5 350.9373743743744u,0 351.9139144144144u,0 351.9149144144144u,1.5 352.8914544544545u,1.5 352.8924544544545u,0 353.8689944944945u,0 353.86999449449445u,1.5 354.8465345345345u,1.5 354.8475345345345u,0 355.8240745745746u,0 355.82507457457456u,1.5 357.7791546546547u,1.5 357.78015465465467u,0 358.7566946946947u,0 358.7576946946947u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 368.5320950950951u,0 368.53309509509506u,1.5 369.50963513513517u,1.5 369.51063513513515u,0 370.4871751751752u,0 370.4881751751752u,1.5 371.4647152152152u,1.5 371.4657152152152u,0 372.44225525525525u,0 372.4432552552552u,1.5 377.3299554554555u,1.5 377.33095545545547u,0 378.3074954954955u,0 378.3084954954955u,1.5 379.28503553553554u,1.5 379.2860355355355u,0 384.1727357357358u,0 384.17373573573576u,1.5 385.15027577577575u,1.5 385.15127577577573u,0 386.1278158158158u,0 386.12881581581576u,1.5 388.0828958958959u,1.5 388.08389589589586u,0 389.06043593593597u,0 389.06143593593595u,1.5 391.99305605605605u,1.5 391.994056056056u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 398.83583633633634u,0 398.8368363363363u,1.5 399.81337637637637u,1.5 399.81437637637634u,0 402.7459964964965u,0 402.7469964964965u,1.5 403.7235365365366u,1.5 403.72453653653656u,0 404.70107657657655u,0 404.70207657657653u,1.5 405.67861661661664u,1.5 405.6796166166166u,0 407.6336966966967u,0 407.63469669669666u,1.5 409.5887767767768u,1.5 409.5897767767768u,0 410.5663168168168u,0 410.5673168168168u,1.5 413.49893693693696u,1.5 413.49993693693693u,0 416.43155705705703u,0 416.432557057057u,1.5 417.40909709709706u,1.5 417.41009709709704u,0 418.38663713713714u,0 418.3876371371371u,1.5 419.36417717717717u,1.5 419.36517717717715u,0 421.3192572572573u,0 421.32025725725725u,1.5 422.29679729729736u,1.5 422.29779729729734u,0 423.27433733733733u,0 423.2753373373373u,1.5 424.25187737737735u,1.5 424.25287737737733u,0 426.20695745745746u,0 426.20795745745744u,1.5 427.18449749749755u,1.5 427.1854974974975u,0 428.16203753753757u,0 428.16303753753755u,1.5 433.04973773773776u,1.5 433.05073773773773u,0 435.98235785785783u,0 435.9833578578578u,1.5 436.9598978978979u,1.5 436.9608978978979u,0 442.82513813813813u,0 442.8261381381381u,1.5 444.78021821821824u,1.5 444.7812182182182u,0 446.73529829829835u,0 446.7362982982983u,1.5 449.6679184184184u,1.5 449.6689184184184u,0 450.64545845845845u,0 450.6464584584584u,1.5 462.37593893893893u,1.5 462.3769389389389u,0 463.353478978979u,0 463.354478978979u,1.5 467.2636391391391u,1.5 467.2646391391391u,0 468.2411791791792u,0 468.2421791791792u,1.5 470.19625925925925u,1.5 470.1972592592592u,0 472.15133933933936u,0 472.15233933933933u,1.5 473.1288793793794u,1.5 473.12987937937936u,0 474.1064194194194u,0 474.1074194194194u,1.5 475.08395945945944u,1.5 475.0849594594594u,0 478.0165795795796u,0 478.0175795795796u,1.5 478.9941196196196u,1.5 478.9951196196196u,0 481.92673973973973u,0 481.9277397397397u,1.5 482.9042797797798u,1.5 482.9052797797798u,0 484.8593598598599u,0 484.8603598598599u,1.5 485.8368998998999u,1.5 485.83789989989987u,0 488.7695200200201u,0 488.77052002002006u,1.5 490.72460010010013u,1.5 490.7256001001001u,0 512.2304809809809u,0 512.2314809809809u,1.5 513.2080210210211u,1.5 513.209021021021u,0 514.1855610610611u,0 514.1865610610611u,1.5 517.1181811811812u,1.5 517.1191811811811u,0 518.0957212212213u,0 518.0967212212213u,1.5 519.0732612612613u,1.5 519.0742612612613u,0 520.0508013013012u,0 520.0518013013012u,1.5 521.0283413413413u,1.5 521.0293413413413u,0 525.9160415415415u,0 525.9170415415415u,1.5 526.8935815815815u,1.5 526.8945815815815u,0 527.8711216216217u,0 527.8721216216217u,1.5 529.8262017017017u,1.5 529.8272017017017u,0 531.7812817817818u,0 531.7822817817818u,1.5 534.7139019019019u,1.5 534.7149019019018u,0 535.6914419419419u,0 535.6924419419419u,1.5 537.646522022022u,1.5 537.647522022022u,0 538.6240620620621u,0 538.625062062062u,1.5 540.5791421421421u,1.5 540.5801421421421u,0 541.5566821821823u,0 541.5576821821822u,1.5 546.4443823823824u,1.5 546.4453823823824u,0 547.4219224224224u,0 547.4229224224224u,1.5 548.3994624624625u,1.5 548.4004624624624u,0 549.3770025025025u,0 549.3780025025025u,1.5 550.3545425425425u,1.5 550.3555425425425u,0 552.3096226226227u,0 552.3106226226226u,1.5 553.2871626626627u,1.5 553.2881626626627u,0 560.1299429429429u,0 560.1309429429429u,1.5 562.085023023023u,1.5 562.086023023023u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 567.9502632632633u,1.5 567.9512632632633u,0 568.9278033033033u,0 568.9288033033033u,1.5 570.8828833833834u,1.5 570.8838833833834u,0 571.8604234234234u,0 571.8614234234234u,1.5 573.8155035035035u,1.5 573.8165035035034u,0 574.7930435435435u,0 574.7940435435435u,1.5 577.7256636636637u,1.5 577.7266636636637u,0 579.6807437437437u,0 579.6817437437437u,1.5 580.6582837837839u,1.5 580.6592837837838u,0 587.501064064064u,0 587.502064064064u,1.5 588.4786041041041u,1.5 588.479604104104u,0 589.4561441441441u,0 589.4571441441441u,1.5 591.4112242242243u,1.5 591.4122242242242u,0 592.3887642642643u,0 592.3897642642643u,1.5 594.3438443443445u,1.5 594.3448443443444u,0 595.3213843843844u,0 595.3223843843843u,1.5 596.2989244244244u,1.5 596.2999244244244u,0 597.2764644644644u,0 597.2774644644644u,1.5 598.2540045045045u,1.5 598.2550045045044u,0 605.0967847847849u,0 605.0977847847848u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 608.0294049049048u,0 608.0304049049048u,1.5 610.962025025025u,1.5 610.963025025025u,0 611.939565065065u,0 611.940565065065u,1.5 613.8946451451452u,1.5 613.8956451451452u,0 614.8721851851852u,0 614.8731851851852u,1.5 615.8497252252253u,1.5 615.8507252252252u,0 619.7598853853854u,0 619.7608853853853u,1.5 620.7374254254254u,1.5 620.7384254254254u,0 621.7149654654654u,0 621.7159654654654u,1.5 622.6925055055054u,1.5 622.6935055055054u,0 623.6700455455456u,0 623.6710455455456u,1.5 626.6026656656657u,1.5 626.6036656656656u,0 627.5802057057057u,0 627.5812057057057u,1.5 629.5352857857858u,1.5 629.5362857857858u,0 633.445445945946u,0 633.4464459459459u,1.5 636.378066066066u,1.5 636.379066066066u,0 637.355606106106u,0 637.356606106106u,1.5 640.2882262262262u,1.5 640.2892262262262u,0 641.2657662662663u,0 641.2667662662662u,1.5 642.2433063063063u,1.5 642.2443063063063u,0 643.2208463463464u,0 643.2218463463464u,1.5 644.1983863863865u,1.5 644.1993863863864u,0 645.1759264264264u,0 645.1769264264263u,1.5 647.1310065065064u,1.5 647.1320065065064u,0 650.0636266266266u,0 650.0646266266266u,1.5 655.9288668668669u,1.5 655.9298668668669u,0 661.7941071071072u,0 661.7951071071071u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 665.7042672672673u,0 665.7052672672672u,1.5 668.6368873873874u,1.5 668.6378873873874u,0 672.5470475475475u,0 672.5480475475475u,1.5 674.5021276276276u,1.5 674.5031276276276u,0 675.4796676676676u,0 675.4806676676676u,1.5 678.4122877877878u,1.5 678.4132877877878u,0 680.3673678678679u,0 680.3683678678678u,1.5 681.344907907908u,1.5 681.345907907908u,0 682.3224479479479u,0 682.3234479479479u,1.5 683.299987987988u,1.5 683.3009879879879u,0 684.277528028028u,0 684.278528028028u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 689.1652282282282u,1.5 689.1662282282282u,0 690.1427682682682u,0 690.1437682682682u,1.5 691.1203083083084u,1.5 691.1213083083084u,0 693.0753883883884u,0 693.0763883883884u,1.5 694.0529284284285u,1.5 694.0539284284284u,0 696.9855485485485u,0 696.9865485485485u,1.5 697.9630885885886u,1.5 697.9640885885885u,0 698.9406286286286u,0 698.9416286286286u,1.5 701.8732487487488u,1.5 701.8742487487488u,0 703.8283288288288u,0 703.8293288288288u,1.5 705.783408908909u,1.5 705.784408908909u,0 709.693569069069u,0 709.694569069069u,1.5 713.6037292292292u,1.5 713.6047292292292u,0 715.5588093093094u,0 715.5598093093093u,1.5 716.5363493493494u,1.5 716.5373493493494u,0 718.4914294294294u,0 718.4924294294294u,1.5 719.4689694694696u,1.5 719.4699694694696u,0 720.4465095095095u,0 720.4475095095095u,1.5 723.3791296296296u,1.5 723.3801296296296u,0 725.3342097097097u,0 725.3352097097097u,1.5 726.3117497497498u,1.5 726.3127497497497u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 730.22190990991u,0 730.22290990991u,1.5 733.15453003003u,1.5 733.1555300300299u,0 734.1320700700701u,0 734.1330700700701u,1.5 736.0871501501501u,1.5 736.0881501501501u,0 739.0197702702703u,0 739.0207702702703u,1.5 743.9074704704706u,1.5 743.9084704704705u,0 745.8625505505505u,0 745.8635505505505u,1.5 746.8400905905905u,1.5 746.8410905905905u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 754.660410910911u,1.5 754.661410910911u,0 755.637950950951u,0 755.638950950951u,1.5 756.615490990991u,1.5 756.616490990991u,0 757.593031031031u,0 757.594031031031u,1.5 759.5481111111111u,1.5 759.5491111111111u,0 761.5031911911911u,0 761.5041911911911u,1.5 763.4582712712713u,1.5 763.4592712712713u,0 766.3908913913914u,0 766.3918913913914u,1.5 767.3684314314314u,1.5 767.3694314314314u,0 768.3459714714716u,0 768.3469714714715u,1.5 769.3235115115116u,1.5 769.3245115115116u,0 770.3010515515515u,0 770.3020515515515u,1.5 774.2112117117117u,1.5 774.2122117117117u,0 775.1887517517517u,0 775.1897517517517u,1.5 776.1662917917918u,1.5 776.1672917917917u,0 778.1213718718719u,0 778.1223718718719u,1.5 779.098911911912u,1.5 779.0999119119119u,0 780.076451951952u,0 780.077451951952u,1.5 781.053991991992u,1.5 781.054991991992u,0 783.0090720720721u,0 783.010072072072u,1.5 785.9416921921921u,1.5 785.9426921921921u,0 786.9192322322323u,0 786.9202322322323u,1.5 787.8967722722723u,1.5 787.8977722722723u,0 791.8069324324325u,0 791.8079324324325u,1.5 796.6946326326326u,1.5 796.6956326326326u,0 797.6721726726727u,0 797.6731726726726u,1.5 798.6497127127127u,1.5 798.6507127127127u,0 799.6272527527527u,0 799.6282527527527u,1.5 800.6047927927928u,1.5 800.6057927927927u,0 801.5823328328329u,0 801.5833328328329u,1.5 802.5598728728729u,1.5 802.5608728728729u,0 803.5374129129129u,0 803.5384129129129u,1.5 804.514952952953u,1.5 804.515952952953u,0 806.4700330330331u,0 806.4710330330331u,1.5 808.4251131131131u,1.5 808.426113113113u,0 811.3577332332333u,0 811.3587332332332u,1.5 812.3352732732733u,1.5 812.3362732732733u,0 813.3128133133133u,0 813.3138133133133u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 816.2454334334335u,0 816.2464334334335u,1.5 817.2229734734735u,1.5 817.2239734734735u,0 818.2005135135136u,0 818.2015135135135u,1.5 820.1555935935936u,1.5 820.1565935935936u,0 822.1106736736737u,0 822.1116736736736u,1.5 823.0882137137137u,1.5 823.0892137137137u,0 825.0432937937937u,0 825.0442937937937u,1.5 826.0208338338339u,1.5 826.0218338338339u,0 826.9983738738739u,0 826.9993738738739u,1.5 830.9085340340341u,1.5 830.9095340340341u,0 832.8636141141141u,0 832.864614114114u,1.5 833.8411541541541u,1.5 833.8421541541541u,0 834.8186941941941u,0 834.8196941941941u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 844.5940945945947u,1.5 844.5950945945947u,0 849.4817947947948u,0 849.4827947947948u,1.5 850.4593348348349u,1.5 850.4603348348348u,0 851.4368748748749u,0 851.4378748748749u,1.5 853.3919549549549u,1.5 853.3929549549549u,0 855.3470350350351u,0 855.3480350350351u,1.5 859.2571951951952u,1.5 859.2581951951952u,0 861.2122752752753u,0 861.2132752752752u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 866.0999754754755u,0 866.1009754754755u,1.5 869.0325955955957u,1.5 869.0335955955957u,0 871.9652157157157u,0 871.9662157157156u,1.5 872.9427557557557u,1.5 872.9437557557557u,0 873.9202957957958u,0 873.9212957957958u,1.5 875.8753758758759u,1.5 875.8763758758759u,0 877.8304559559559u,0 877.8314559559559u,1.5 878.8079959959961u,1.5 878.808995995996u,0 879.7855360360361u,0 879.7865360360361u,1.5 885.6507762762762u,1.5 885.6517762762762u,0 886.6283163163163u,0 886.6293163163162u,1.5 887.6058563563563u,1.5 887.6068563563563u,0 895.4261766766766u,0 895.4271766766766u,1.5 898.3587967967968u,1.5 898.3597967967968u,0 899.3363368368368u,0 899.3373368368368u,1.5 900.3138768768769u,1.5 900.3148768768768u,0 901.2914169169169u,0 901.2924169169169u,1.5 902.2689569569569u,1.5 902.2699569569569u,0 903.246496996997u,0 903.247496996997u,1.5 904.2240370370371u,1.5 904.225037037037u,0 905.2015770770771u,0 905.2025770770771u,1.5 907.1566571571572u,1.5 907.1576571571571u,0 910.0892772772772u,0 910.0902772772772u,1.5 913.9994374374375u,1.5 914.0004374374374u,0 915.9545175175175u,0 915.9555175175175u,1.5 918.8871376376377u,1.5 918.8881376376377u,0 919.8646776776777u,0 919.8656776776777u,1.5 920.8422177177176u,1.5 920.8432177177176u,0 921.8197577577578u,0 921.8207577577577u,1.5 922.7972977977978u,1.5 922.7982977977978u,0 928.6625380380381u,0 928.663538038038u,1.5 930.6176181181181u,1.5 930.6186181181181u,0 934.5277782782782u,0 934.5287782782782u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 936.4828583583584u,0 936.4838583583584u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 940.3930185185185u,0 940.3940185185185u,1.5 946.2582587587588u,1.5 946.2592587587587u,0 947.2357987987988u,0 947.2367987987988u,1.5 948.2133388388388u,1.5 948.2143388388388u,0 950.1684189189189u,0 950.1694189189188u,1.5 951.145958958959u,1.5 951.146958958959u,0 952.123498998999u,0 952.124498998999u,1.5 953.101039039039u,1.5 953.102039039039u,0 954.0785790790791u,0 954.079579079079u,1.5 955.0561191191191u,1.5 955.0571191191191u,0 960.9213593593594u,0 960.9223593593593u,1.5 962.8764394394394u,1.5 962.8774394394394u,0 964.8315195195195u,0 964.8325195195195u,1.5 965.8090595595596u,1.5 965.8100595595596u,0 968.7416796796797u,0 968.7426796796797u,1.5 970.6967597597597u,1.5 970.6977597597597u,0 972.6518398398398u,0 972.6528398398398u,1.5 973.6293798798798u,1.5 973.6303798798798u,0 974.60691991992u,0 974.6079199199199u,1.5 975.58445995996u,1.5 975.58545995996u,0 976.562u,0 976.563u,1.5 977.5395400400402u,1.5 977.5405400400401u,0 978.5170800800801u,0 978.51808008008u,1.5 982.4272402402403u,1.5 982.4282402402403u,0 983.4047802802802u,0 983.4057802802802u,1.5 984.3823203203203u,1.5 984.3833203203203u,0 985.3598603603602u,0 985.3608603603602u,1.5 986.3374004004004u,1.5 986.3384004004004u,0 987.3149404404405u,0 987.3159404404405u,1.5 988.2924804804804u,1.5 988.2934804804804u,0 989.2700205205206u,0 989.2710205205206u,1.5 993.1801806806807u,1.5 993.1811806806807u,0 994.1577207207208u,0 994.1587207207208u,1.5 997.0903408408409u,1.5 997.0913408408409u,0 998.0678808808808u,0 998.0688808808808u,1.5 999.045420920921u,1.5 999.0464209209209u,0 1001.9780410410411u,0 1001.9790410410411u,1.5 1011.7534414414415u,1.5 1011.7544414414415u,0 1014.6860615615615u,0 1014.6870615615614u,1.5 1021.5288418418419u,1.5 1021.5298418418419u,0 1022.5063818818818u,0 1022.5073818818818u,1.5 1023.4839219219219u,1.5 1023.4849219219219u,0 1025.4390020020019u,0 1025.440002002002u,1.5 1026.416542042042u,1.5 1026.4175420420422u,0 1027.394082082082u,0 1027.3950820820821u,1.5 1028.371622122122u,1.5 1028.3726221221223u,0 1029.349162162162u,0 1029.3501621621622u,1.5 1030.3267022022021u,1.5 1030.3277022022023u,0 1031.3042422422423u,0 1031.3052422422425u,1.5 1032.2817822822822u,1.5 1032.2827822822824u,0 1034.2368623623622u,0 1034.2378623623624u,1.5 1035.2144024024024u,1.5 1035.2154024024026u,0 1038.1470225225225u,0 1038.1480225225228u,1.5 1039.1245625625625u,1.5 1039.1255625625627u,0 1042.0571826826824u,0 1042.0581826826826u,1.5 1043.0347227227226u,1.5 1043.0357227227228u,0 1045.9673428428428u,0 1045.968342842843u,1.5 1046.9448828828827u,1.5 1046.9458828828829u,0 1047.9224229229228u,0 1047.923422922923u,1.5 1048.8999629629627u,1.5 1048.900962962963u,0 1049.8775030030029u,0 1049.878503003003u,1.5 1050.855043043043u,1.5 1050.8560430430432u,0 1051.832583083083u,0 1051.833583083083u,1.5 1052.810123123123u,1.5 1052.8111231231233u,0 1053.787663163163u,0 1053.7886631631632u,1.5 1055.7427432432432u,1.5 1055.7437432432434u,0 1056.7202832832832u,0 1056.7212832832834u,1.5 1063.5630635635634u,1.5 1063.5640635635636u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1073.338463963964u,0 1073.3394639639641u,1.5 1074.3160040040038u,1.5 1074.317004004004u,0 1077.248624124124u,0 1077.2496241241242u,1.5 1085.0689444444445u,1.5 1085.0699444444447u,0 1088.9791046046046u,0 1088.9801046046048u,1.5 1089.9566446446445u,1.5 1089.9576446446447u,0 1091.9117247247245u,0 1091.9127247247247u,1.5 1092.8892647647647u,1.5 1092.8902647647649u,0 1093.8668048048046u,0 1093.8678048048048u,1.5 1095.8218848848846u,1.5 1095.8228848848848u,0 1096.7994249249248u,0 1096.800424924925u,1.5 1099.732045045045u,1.5 1099.7330450450452u,0 1100.7095850850849u,0 1100.710585085085u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1112.4400655655656u,0 1112.4410655655659u,1.5 1113.4176056056056u,1.5 1113.4186056056058u,0 1115.3726856856854u,0 1115.3736856856856u,1.5 1120.2603858858856u,1.5 1120.2613858858858u,0 1121.2379259259258u,0 1121.238925925926u,1.5 1122.215465965966u,1.5 1122.216465965966u,0 1123.1930060060058u,0 1123.194006006006u,1.5 1124.170546046046u,1.5 1124.1715460460462u,0 1126.125626126126u,0 1126.1266261261262u,1.5 1128.080706206206u,1.5 1128.0817062062063u,0 1130.035786286286u,0 1130.0367862862863u,1.5 1131.0133263263263u,1.5 1131.0143263263265u,0 1131.9908663663664u,0 1131.9918663663666u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1137.8561066066065u,1.5 1137.8571066066067u,0 1140.7887267267265u,0 1140.7897267267267u,1.5 1141.7662667667666u,1.5 1141.7672667667669u,0 1143.7213468468467u,0 1143.722346846847u,1.5 1145.6764269269268u,1.5 1145.677426926927u,0 1146.653966966967u,0 1146.654966966967u,1.5 1148.609047047047u,1.5 1148.6100470470471u,0 1149.5865870870869u,0 1149.587587087087u,1.5 1150.564127127127u,1.5 1150.5651271271272u,0 1156.4293673673674u,0 1156.4303673673676u,1.5 1157.4069074074073u,1.5 1157.4079074074075u,0 1158.3844474474474u,0 1158.3854474474476u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1169.1373878878876u,0 1169.1383878878878u,1.5 1174.0250880880878u,1.5 1174.026088088088u,0 1175.9801681681681u,0 1175.9811681681683u,1.5 1176.957708208208u,1.5 1176.9587082082082u,0 1177.9352482482482u,0 1177.9362482482484u,1.5 1178.912788288288u,1.5 1178.9137882882883u,0 1179.8903283283282u,0 1179.8913283283284u,1.5 1180.8678683683684u,1.5 1180.8688683683686u,0 1183.8004884884883u,0 1183.8014884884885u,1.5 1184.7780285285285u,1.5 1184.7790285285287u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1186.7331086086085u,1.5 1186.7341086086087u,0 1191.6208088088085u,0 1191.6218088088087u,1.5 1193.5758888888888u,1.5 1193.576888888889u,0 1194.5534289289287u,0 1194.554428928929u,1.5 1195.5309689689689u,1.5 1195.531968968969u,0 1196.5085090090088u,0 1196.509509009009u,1.5 1197.486049049049u,1.5 1197.4870490490491u,0 1201.396209209209u,0 1201.3972092092092u,1.5 1202.3737492492492u,1.5 1202.3747492492494u,0 1203.3512892892893u,0 1203.3522892892895u,1.5 1204.3288293293292u,1.5 1204.3298293293294u,0 1205.3063693693693u,0 1205.3073693693696u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1212.1491496496496u,0 1212.1501496496498u,1.5 1213.1266896896898u,1.5 1213.12768968969u,0 1216.0593098098095u,0 1216.0603098098097u,1.5 1217.0368498498497u,1.5 1217.0378498498499u,0 1218.0143898898898u,0 1218.01538988989u,1.5 1218.9919299299297u,1.5 1218.99292992993u,0 1222.90209009009u,0 1222.9030900900902u,1.5 1223.87963013013u,1.5 1223.8806301301302u,0 1225.83471021021u,0 1225.8357102102102u,1.5 1227.7897902902903u,1.5 1227.7907902902905u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1234.6325705705706u,0 1234.6335705705708u,1.5 1239.5202707707706u,1.5 1239.5212707707708u,0 1241.4753508508506u,0 1241.4763508508508u,1.5 1242.4528908908908u,1.5 1242.453890890891u,0 1245.3855110110107u,0 1245.386511011011u,1.5 1247.340591091091u,1.5 1247.3415910910912u,0 1248.318131131131u,0 1248.3191311311311u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1256.1384514514514u,0 1256.1394514514516u,1.5 1259.0710715715716u,1.5 1259.0720715715718u,0 1261.0261516516516u,0 1261.0271516516518u,1.5 1262.0036916916918u,1.5 1262.004691691692u,0 1262.9812317317317u,0 1262.9822317317319u,1.5 1263.9587717717718u,1.5 1263.959771771772u,0 1264.9363118118117u,0 1264.937311811812u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1269.8240120120117u,0 1269.825012012012u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1274.711712212212u,0 1274.7127122122122u,1.5 1275.6892522522521u,1.5 1275.6902522522523u,0 1276.6667922922923u,0 1276.6677922922925u,1.5 1282.5320325325324u,1.5 1282.5330325325326u,0 1287.4197327327327u,0 1287.4207327327329u,1.5 1288.3972727727728u,1.5 1288.398272772773u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1296.217593093093u,1.5 1296.2185930930932u,0 1297.195133133133u,0 1297.1961331331331u,1.5 1298.172673173173u,1.5 1298.1736731731733u,0 1300.127753253253u,0 1300.1287532532533u,1.5 1301.1052932932932u,1.5 1301.1062932932934u,0 1302.0828333333332u,0 1302.0838333333334u,1.5 1303.0603733733733u,1.5 1303.0613733733735u,0 1305.0154534534533u,0 1305.0164534534536u,1.5 1306.9705335335334u,1.5 1306.9715335335336u,0 1308.9256136136135u,0 1308.9266136136137u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1320.656094094094u,0 1320.6570940940942u,1.5 1321.633634134134u,1.5 1321.634634134134u,0 1322.611174174174u,0 1322.6121741741742u,1.5 1324.566254254254u,1.5 1324.5672542542543u,0 1325.5437942942942u,0 1325.5447942942944u,1.5 1326.5213343343341u,1.5 1326.5223343343343u,0 1332.3865745745745u,0 1332.3875745745747u,1.5 1336.2967347347346u,1.5 1336.2977347347348u,0 1337.2742747747748u,0 1337.275274774775u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1340.2068948948947u,0 1340.207894894895u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1344.1170550550548u,0 1344.118055055055u,1.5 1345.094595095095u,1.5 1345.0955950950952u,0 1346.0721351351349u,0 1346.073135135135u,1.5 1350.9598353353351u,1.5 1350.9608353353353u,0 1352.9149154154154u,0 1352.9159154154156u,1.5 1353.8924554554553u,1.5 1353.8934554554555u,0 1354.8699954954955u,0 1354.8709954954957u,1.5 1355.8475355355354u,1.5 1355.8485355355356u,0 1356.8250755755755u,0 1356.8260755755757u,1.5 1358.7801556556556u,1.5 1358.7811556556558u,0 1359.7576956956957u,0 1359.758695695696u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1363.6678558558558u,1.5 1363.668855855856u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1365.6229359359356u,1.5 1365.6239359359358u,0 1370.5106361361359u,0 1370.511636136136u,1.5 1371.488176176176u,1.5 1371.4891761761762u,0 1372.4657162162162u,0 1372.4667162162164u,1.5 1378.3309564564563u,1.5 1378.3319564564565u,0 1380.2860365365364u,0 1380.2870365365366u,1.5 1381.2635765765765u,1.5 1381.2645765765767u,0 1383.2186566566565u,0 1383.2196566566568u,1.5 1384.1961966966967u,1.5 1384.197196696697u,0 1385.1737367367366u,0 1385.1747367367368u,1.5 1387.1288168168169u,1.5 1387.129816816817u,0 1388.1063568568568u,0 1388.107356856857u,1.5 1391.0389769769768u,1.5 1391.039976976977u,0 1392.016517017017u,0 1392.017517017017u,1.5 1392.9940570570568u,1.5 1392.995057057057u,0 1393.971597097097u,0 1393.9725970970972u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1395.926677177177u,0 1395.9276771771772u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1401.7919174174174u,0 1401.7929174174176u,1.5 1403.7469974974974u,1.5 1403.7479974974976u,0 1405.7020775775775u,0 1405.7030775775777u,1.5 1408.6346976976977u,1.5 1408.6356976976979u,0 1409.6122377377376u,0 1409.6132377377378u,1.5 1412.5448578578578u,1.5 1412.545857857858u,0 1413.522397897898u,0 1413.5233978978981u,1.5 1415.4774779779777u,1.5 1415.478477977978u,0 1416.4550180180179u,0 1416.456018018018u,1.5 1419.3876381381378u,1.5 1419.388638138138u,0 1420.365178178178u,0 1420.3661781781782u,1.5 1422.320258258258u,1.5 1422.3212582582582u,0 1423.2977982982982u,0 1423.2987982982984u,1.5 1424.275338338338u,1.5 1424.2763383383383u,0 1425.2528783783782u,0 1425.2538783783784u,1.5 1436.9833588588588u,1.5 1436.984358858859u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1440.8935190190189u,1.5 1440.894519019019u,0 1441.8710590590588u,0 1441.872059059059u,1.5 1443.826139139139u,1.5 1443.8271391391393u,0 1447.7362992992992u,0 1447.7372992992994u,1.5 1453.6015395395395u,1.5 1453.6025395395397u,0 1454.5790795795795u,0 1454.5800795795797u,1.5 1463.37693993994u,1.5 1463.3779399399402u,0 1464.35447997998u,0 1464.3554799799801u,1.5 1466.3095600600598u,1.5 1466.31056006006u,0 1467.2871001001u,0 1467.2881001001u,1.5 1468.26464014014u,1.5 1468.2656401401402u,0 1469.24218018018u,0 1469.2431801801802u,1.5 1476.0849604604603u,1.5 1476.0859604604605u,0 1478.0400405405405u,0 1478.0410405405407u,1.5 1479.0175805805804u,1.5 1479.0185805805806u,0 1482.9277407407408u,0 1482.928740740741u,1.5 1483.9052807807807u,1.5 1483.906280780781u,0 1486.8379009009009u,0 1486.838900900901u,1.5 1487.815440940941u,1.5 1487.8164409409412u,0 1488.792980980981u,0 1488.7939809809811u,1.5 1489.7705210210208u,1.5 1489.771521021021u,0 1493.680681181181u,0 1493.6816811811811u,1.5 1495.635761261261u,1.5 1495.6367612612612u,0 1496.6133013013011u,0 1496.6143013013013u,1.5 1498.5683813813812u,1.5 1498.5693813813814u,0 1499.5459214214213u,0 1499.5469214214215u,1.5 1500.5234614614612u,1.5 1500.5244614614614u,0 1501.5010015015014u,0 1501.5020015015016u,1.5 1502.4785415415415u,1.5 1502.4795415415417u,0 1506.3887017017016u,0 1506.3897017017018u,1.5 1508.3437817817817u,1.5 1508.3447817817819u,0 1512.253941941942u,0 1512.2549419419422u,1.5 1513.231481981982u,1.5 1513.2324819819821u,0 1514.209022022022u,0 1514.2100220220223u,1.5 1515.186562062062u,1.5 1515.1875620620622u,0 1521.0518023023021u,0 1521.0528023023023u,1.5 1522.0293423423423u,1.5 1522.0303423423425u,0 1525.9395025025024u,0 1525.9405025025026u,1.5 1528.8721226226226u,1.5 1528.8731226226228u,0 1529.8496626626625u,0 1529.8506626626627u,1.5 1530.8272027027026u,1.5 1530.8282027027028u,0 1531.8047427427427u,0 1531.805742742743u,1.5 1534.7373628628627u,1.5 1534.738362862863u,0 1535.7149029029028u,0 1535.715902902903u,1.5 1537.669982982983u,1.5 1537.670982982983u,0 1538.647523023023u,0 1538.6485230230232u,1.5 1539.625063063063u,1.5 1539.6260630630632u,0 1542.557683183183u,0 1542.5586831831831u,1.5 1546.4678433433432u,1.5 1546.4688433433435u,0 1547.4453833833832u,0 1547.4463833833834u,1.5 1549.4004634634632u,1.5 1549.4014634634634u,0 1550.3780035035034u,0 1550.3790035035036u,1.5 1551.3555435435435u,1.5 1551.3565435435437u,0 1552.3330835835834u,0 1552.3340835835836u,1.5 1553.3106236236235u,1.5 1553.3116236236237u,0 1556.2432437437437u,0 1556.244243743744u,1.5 1557.2207837837836u,1.5 1557.2217837837838u,0 1561.130943943944u,0 1561.1319439439442u,1.5 1563.086024024024u,1.5 1563.0870240240242u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1566.018644144144u,1.5 1566.0196441441442u,0 1566.996184184184u,0 1566.997184184184u,1.5 1577.7491246246245u,1.5 1577.7501246246247u,0 1581.6592847847846u,0 1581.6602847847848u,1.5 1582.6368248248248u,1.5 1582.637824824825u,0 1583.614364864865u,0 1583.6153648648651u,1.5 1584.5919049049048u,1.5 1584.592904904905u,0 1587.524525025025u,0 1587.5255250250252u,1.5 1589.479605105105u,1.5 1589.4806051051053u,0 1590.457145145145u,0 1590.4581451451452u,1.5 1596.3223853853851u,1.5 1596.3233853853853u,0 1598.2774654654654u,0 1598.2784654654656u,1.5 1599.2550055055053u,1.5 1599.2560055055055u,0 1600.2325455455455u,0 1600.2335455455457u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1610.9854859859859u,1.5 1610.986485985986u,0 1611.963026026026u,0 1611.9640260260262u,1.5 1612.9405660660661u,1.5 1612.9415660660663u,0 1614.8956461461462u,0 1614.8966461461464u,1.5 1615.8731861861859u,1.5 1615.874186186186u,0 1616.850726226226u,0 1616.8517262262262u,1.5 1617.8282662662662u,1.5 1617.8292662662664u,0 1619.7833463463462u,0 1619.7843463463464u,1.5 1620.7608863863861u,1.5 1620.7618863863863u,0 1621.7384264264263u,0 1621.7394264264265u,1.5 1622.7159664664664u,1.5 1622.7169664664666u,0 1623.6935065065063u,0 1623.6945065065065u,1.5 1624.6710465465464u,1.5 1624.6720465465467u,0 1625.6485865865864u,0 1625.6495865865866u,1.5 1628.5812067067066u,1.5 1628.5822067067068u,0 1629.5587467467467u,0 1629.559746746747u,1.5 1630.5362867867866u,1.5 1630.5372867867868u,0 1633.4689069069068u,0 1633.469906906907u,1.5 1634.446446946947u,1.5 1634.4474469469471u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1639.3341471471472u,1.5 1639.3351471471474u,0 1640.311687187187u,0 1640.3126871871873u,1.5 1642.2667672672671u,1.5 1642.2677672672673u,0 1644.2218473473472u,0 1644.2228473473474u,1.5 1645.199387387387u,1.5 1645.2003873873873u,0 1649.1095475475474u,0 1649.1105475475476u,1.5 1651.0646276276275u,1.5 1651.0656276276277u,0 1652.0421676676676u,0 1652.0431676676678u,1.5 1655.9523278278277u,1.5 1655.953327827828u,0 1656.9298678678679u,0 1656.930867867868u,1.5 1657.9074079079078u,1.5 1657.908407907908u,0 1658.884947947948u,0 1658.8859479479481u,1.5 1660.840028028028u,1.5 1660.8410280280282u,0 1664.750188188188u,0 1664.7511881881883u,1.5 1667.682808308308u,1.5 1667.6838083083082u,0 1674.5255885885883u,0 1674.5265885885885u,1.5 1680.3908288288287u,1.5 1680.391828828829u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1686.256069069069u,1.5 1686.2570690690693u,0 1687.233609109109u,0 1687.2346091091092u,1.5 1691.1437692692691u,1.5 1691.1447692692693u,0 1696.0314694694694u,0 1696.0324694694696u,1.5 1697.9865495495494u,1.5 1697.9875495495496u,0 1698.9640895895895u,0 1698.9650895895898u,1.5 1701.8967097097095u,1.5 1701.8977097097097u,0 1702.8742497497497u,0 1702.8752497497499u,1.5 1703.8517897897898u,1.5 1703.85278978979u,0 1704.8293298298297u,0 1704.83032982983u,1.5 1705.8068698698698u,1.5 1705.80786986987u,0 1706.7844099099098u,0 1706.78540990991u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1708.73948998999u,0 1708.7404899899902u,1.5 1710.69457007007u,1.5 1710.6955700700703u,0 1717.5373503503502u,0 1717.5383503503504u,1.5 1718.5148903903903u,1.5 1718.5158903903905u,0 1719.4924304304302u,0 1719.4934304304304u,1.5 1727.3127507507506u,1.5 1727.3137507507508u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1731.2229109109107u,1.5 1731.223910910911u,0 1732.2004509509509u,0 1732.201450950951u,1.5 1733.177990990991u,1.5 1733.1789909909912u,0 1739.0432312312312u,0 1739.0442312312314u,1.5 1740.0207712712713u,1.5 1740.0217712712715u,0 1740.998311311311u,0 1740.9993113113112u,1.5 1741.9758513513511u,1.5 1741.9768513513513u,0 1743.9309314314312u,0 1743.9319314314314u,1.5 1745.8860115115112u,1.5 1745.8870115115114u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1755.6614119119117u,1.5 1755.662411911912u,0 1760.549112112112u,0 1760.5501121121122u,1.5 1762.5041921921922u,1.5 1762.5051921921925u,0 1763.4817322322322u,0 1763.4827322322324u,1.5 1765.4368123123122u,1.5 1765.4378123123124u,0 1770.3245125125122u,0 1770.3255125125124u,1.5 1772.2795925925925u,1.5 1772.2805925925927u,0 1773.2571326326324u,0 1773.2581326326326u,1.5 1774.2346726726726u,1.5 1774.2356726726728u,0 1776.1897527527526u,0 1776.1907527527528u,1.5 1777.1672927927928u,1.5 1777.168292792793u,0 1778.1448328328327u,0 1778.1458328328329u,1.5 1779.1223728728728u,1.5 1779.123372872873u,0 1782.054992992993u,0 1782.0559929929932u,1.5 1787.9202332332331u,1.5 1787.9212332332334u,0 1788.8977732732733u,0 1788.8987732732735u,1.5 1789.8753133133132u,1.5 1789.8763133133134u,0 1791.8303933933933u,0 1791.8313933933935u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1797.6956336336334u,1.5 1797.6966336336336u,0 1798.6731736736735u,0 1798.6741736736737u,1.5 1799.6507137137135u,1.5 1799.6517137137137u,0 1800.6282537537536u,0 1800.6292537537538u,1.5 1801.6057937937937u,1.5 1801.606793793794u,0 1804.5384139139137u,0 1804.539413913914u,1.5 1806.493493993994u,1.5 1806.4944939939942u,0 1807.471034034034u,0 1807.472034034034u,1.5 1808.448574074074u,1.5 1808.4495740740742u,0 1809.426114114114u,0 1809.4271141141141u,1.5 1810.403654154154u,1.5 1810.4046541541543u,0 1811.3811941941942u,0 1811.3821941941944u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1814.3138143143142u,1.5 1814.3148143143144u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1820.1790545545543u,1.5 1820.1800545545545u,0 1821.1565945945945u,0 1821.1575945945947u,1.5 1822.1341346346344u,1.5 1822.1351346346346u,0 1823.1116746746745u,0 1823.1126746746747u,1.5 1824.0892147147147u,1.5 1824.0902147147149u,0 1826.0442947947947u,0 1826.045294794795u,1.5 1827.9993748748748u,1.5 1828.000374874875u,0 1829.9544549549548u,0 1829.955454954955u,1.5 1830.931994994995u,1.5 1830.9329949949952u,0 1831.9095350350349u,0 1831.910535035035u,1.5 1832.887075075075u,1.5 1832.8880750750752u,0 1833.8646151151152u,0 1833.8656151151154u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1843.6400155155154u,1.5 1843.6410155155156u,0 1844.6175555555553u,0 1844.6185555555555u,1.5 1845.5950955955955u,1.5 1845.5960955955957u,0 1851.4603358358356u,0 1851.4613358358358u,1.5 1855.370495995996u,1.5 1855.3714959959962u,0 1857.325576076076u,0 1857.3265760760762u,1.5 1858.3031161161161u,1.5 1858.3041161161163u,0 1859.280656156156u,0 1859.2816561561563u,1.5 1860.2581961961962u,1.5 1860.2591961961964u,0 1861.235736236236u,0 1861.2367362362363u,1.5 1862.2132762762762u,1.5 1862.2142762762765u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1867.1009764764763u,1.5 1867.1019764764765u,0 1868.0785165165164u,0 1868.0795165165166u,1.5 1871.0111366366364u,1.5 1871.0121366366366u,0 1872.9662167167166u,0 1872.9672167167168u,1.5 1873.9437567567566u,1.5 1873.9447567567568u,0 1876.8763768768767u,0 1876.877376876877u,1.5 1877.853916916917u,1.5 1877.854916916917u,0 1878.8314569569568u,0 1878.832456956957u,1.5 1880.7865370370369u,1.5 1880.787537037037u,0 1882.7416171171171u,0 1882.7426171171173u,1.5 1884.6966971971972u,1.5 1884.6976971971974u,0 1885.674237237237u,0 1885.6752372372373u,1.5 1888.6068573573573u,1.5 1888.6078573573575u,0 1889.5843973973974u,0 1889.5853973973976u,1.5 1891.5394774774772u,1.5 1891.5404774774775u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1895.4496376376374u,0 1895.4506376376376u,1.5 1900.3373378378376u,1.5 1900.3383378378378u,0 1901.3148778778777u,0 1901.315877877878u,1.5 1903.2699579579578u,1.5 1903.270957957958u,0 1906.202578078078u,0 1906.2035780780782u,1.5 1907.1801181181181u,1.5 1907.1811181181183u,0 1913.0453583583583u,0 1913.0463583583585u,1.5 1914.0228983983984u,1.5 1914.0238983983986u,0 1915.0004384384383u,0 1915.0014384384385u,1.5 1921.8432187187186u,1.5 1921.8442187187188u,0 1924.7758388388386u,0 1924.7768388388388u,1.5 1925.7533788788787u,1.5 1925.754378878879u,0 1928.685998998999u,0 1928.6869989989991u,1.5 1929.6635390390388u,1.5 1929.664539039039u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1934.551239239239u,0 1934.5522392392393u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1939.4389394394395u,0 1939.4399394394397u,1.5 1942.3715595595593u,1.5 1942.3725595595595u,0 1943.3490995995994u,0 1943.3500995995996u,1.5 1947.2592597597595u,1.5 1947.2602597597597u,0 1948.2367997997997u,0 1948.2377997997999u,1.5 1950.1918798798797u,1.5 1950.19287987988u,0 1951.1694199199198u,0 1951.17041991992u,1.5 1952.1469599599598u,1.5 1952.14795995996u,0 1953.1245u,0 1953.1255u,1.5 1954.10204004004u,1.5 1954.1030400400402u,0 1955.0795800800802u,0 1955.0805800800804u,1.5 1956.0571201201199u,1.5 1956.05812012012u,0 1959.9672802802804u,0 1959.9682802802806u,1.5 1961.9223603603602u,1.5 1961.9233603603604u,0 1967.7876006006004u,0 1967.7886006006006u,1.5 1969.7426806806807u,1.5 1969.7436806806809u,0 1970.7202207207204u,0 1970.7212207207206u,1.5 1971.6977607607605u,1.5 1971.6987607607607u,0 1972.6753008008006u,0 1972.6763008008008u,1.5 1973.6528408408408u,1.5 1973.653840840841u,0 1974.630380880881u,0 1974.6313808808811u,1.5 1975.6079209209206u,1.5 1975.6089209209208u,0 1976.5854609609607u,0 1976.586460960961u,1.5 1978.540541041041u,1.5 1978.5415410410412u,0 1979.5180810810812u,0 1979.5190810810814u,1.5 1982.4507012012011u,1.5 1982.4517012012013u,0 1983.4282412412413u,0 1983.4292412412415u,1.5 1988.3159414414415u,1.5 1988.3169414414417u,0 1989.2934814814816u,0 1989.2944814814819u,1.5 1995.1587217217213u,1.5 1995.1597217217216u,0 1996.1362617617615u,0 1996.1372617617617u,1.5 1997.1138018018016u,1.5 1997.1148018018018u,0 1999.068881881882u,0 1999.069881881882u,1.5 2002.979042042042u,1.5 2002.9800420420422u,0 2003.9565820820822u,0 2003.9575820820824u,1.5 2005.911662162162u,1.5 2005.9126621621622u,0 2006.8892022022021u,0 2006.8902022022023u,1.5 2017.6421426426425u,1.5 2017.6431426426427u,0 2018.6196826826827u,0 2018.6206826826829u,1.5 2020.5747627627625u,1.5 2020.5757627627627u,0 2021.5523028028026u,0 2021.5533028028028u,1.5 2024.4849229229226u,1.5 2024.4859229229228u,0 2025.4624629629627u,0 2025.463462962963u,1.5 2027.417543043043u,1.5 2027.4185430430432u,0 2030.350163163163u,0 2030.3511631631632u,1.5 2031.327703203203u,1.5 2031.3287032032033u,0 2032.3052432432432u,0 2032.3062432432434u,1.5 2033.2827832832834u,1.5 2033.2837832832836u,0 2038.1704834834836u,0 2038.1714834834838u,1.5 2039.1480235235233u,1.5 2039.1490235235235u,0 2045.9908038038036u,0 2045.9918038038038u,1.5 2046.9683438438437u,1.5 2046.969343843844u,0 2049.900963963964u,0 2049.901963963964u,1.5 2050.878504004004u,1.5 2050.879504004004u,0 2053.811124124124u,0 2053.8121241241242u,1.5 2058.698824324324u,1.5 2058.6998243243243u,0 2059.676364364364u,0 2059.677364364364u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2065.5416046046043u,0 2065.5426046046045u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2069.4517647647644u,1.5 2069.4527647647647u,0 2072.384384884885u,0 2072.3853848848853u,1.5 2074.339464964965u,1.5 2074.340464964965u,0 2076.294545045045u,0 2076.2955450450454u,1.5 2077.272085085085u,1.5 2077.2730850850853u,0 2078.249625125125u,0 2078.250625125125u,1.5 2088.025025525525u,1.5 2088.0260255255253u,0 2095.8453458458457u,0 2095.846345845846u,1.5 2097.8004259259255u,1.5 2097.8014259259257u,0 2098.777965965966u,0 2098.778965965966u,1.5 2099.755506006006u,1.5 2099.756506006006u,0 2100.733046046046u,0 2100.7340460460464u,1.5 2103.665666166166u,1.5 2103.666666166166u,0 2107.575826326326u,0 2107.576826326326u,1.5 2108.553366366366u,1.5 2108.554366366366u,0 2111.4859864864866u,0 2111.486986486487u,1.5 2115.3961466466467u,1.5 2115.397146646647u,0 2117.3512267267265u,0 2117.3522267267267u,1.5 2122.2389269269265u,1.5 2122.2399269269267u,0 2123.216466966967u,0 2123.217466966967u,1.5 2127.126627127127u,1.5 2127.127627127127u,0 2128.104167167167u,0 2128.105167167167u,1.5 2129.081707207207u,1.5 2129.082707207207u,0 2130.059247247247u,0 2130.0602472472474u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2138.8571076076073u,0 2138.8581076076075u,1.5 2139.8346476476477u,1.5 2139.835647647648u,0 2142.7672677677674u,0 2142.7682677677676u,1.5 2143.744807807808u,1.5 2143.745807807808u,0 2144.7223478478477u,0 2144.723347847848u,1.5 2147.654967967968u,1.5 2147.655967967968u,0 2148.632508008008u,0 2148.633508008008u,1.5 2149.610048048048u,1.5 2149.6110480480484u,0 2156.4528283283285u,0 2156.4538283283287u,1.5 2157.430368368368u,1.5 2157.431368368368u,0 2158.4079084084083u,0 2158.4089084084085u,1.5 2159.385448448448u,1.5 2159.3864484484484u,0 2160.3629884884886u,0 2160.3639884884888u,1.5 2161.3405285285285u,1.5 2161.3415285285287u,0 2166.228228728729u,0 2166.229228728729u,1.5 2168.1833088088088u,1.5 2168.184308808809u,0 2169.1608488488487u,0 2169.161848848849u,1.5 2171.115928928929u,1.5 2171.116928928929u,0 2173.071009009009u,0 2173.072009009009u,1.5 2175.026089089089u,1.5 2175.0270890890893u,0 2177.9587092092092u,0 2177.9597092092094u,1.5 2178.936249249249u,1.5 2178.9372492492494u,0 2179.913789289289u,0 2179.9147892892893u,1.5 2180.8913293293294u,1.5 2180.8923293293296u,0 2181.868869369369u,0 2181.869869369369u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2189.6891896896896u,0 2189.6901896896898u,1.5 2190.66672972973u,1.5 2190.66772972973u,0 2191.6442697697694u,0 2191.6452697697696u,1.5 2196.53196996997u,1.5 2196.53296996997u,0 2198.48705005005u,0 2198.4880500500503u,1.5 2199.46459009009u,1.5 2199.4655900900902u,0 2200.4421301301304u,0 2200.4431301301306u,1.5 2203.37475025025u,1.5 2203.3757502502503u,0 2204.35229029029u,0 2204.3532902902903u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2211.1950705705704u,0 2211.1960705705706u,1.5 2212.1726106106103u,1.5 2212.1736106106105u,0 2213.1501506506506u,0 2213.151150650651u,1.5 2215.105230730731u,1.5 2215.106230730731u,0 2216.0827707707704u,0 2216.0837707707706u,1.5 2219.015390890891u,1.5 2219.016390890891u,0 2222.925551051051u,0 2222.9265510510513u,1.5 2223.903091091091u,1.5 2223.9040910910912u,0 2224.8806311311314u,0 2224.8816311311316u,1.5 2225.858171171171u,1.5 2225.859171171171u,0 2226.835711211211u,0 2226.8367112112114u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2232.700951451451u,0 2232.7019514514514u,1.5 2242.4763518518516u,1.5 2242.477351851852u,0 2244.431431931932u,0 2244.432431931932u,1.5 2245.408971971972u,1.5 2245.409971971972u,0 2246.3865120120117u,0 2246.387512012012u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2255.184372372372u,0 2255.185372372372u,1.5 2256.161912412412u,1.5 2256.1629124124124u,0 2257.139452452452u,0 2257.1404524524523u,1.5 2258.1169924924925u,1.5 2258.1179924924927u,0 2259.0945325325324u,0 2259.0955325325326u,1.5 2261.0496126126122u,1.5 2261.0506126126124u,0 2262.0271526526526u,0 2262.028152652653u,1.5 2263.0046926926925u,1.5 2263.0056926926927u,0 2263.982232732733u,0 2263.983232732733u,1.5 2264.9597727727723u,1.5 2264.9607727727725u,0 2265.9373128128127u,0 2265.938312812813u,1.5 2266.9148528528526u,1.5 2266.915852852853u,0 2267.892392892893u,0 2267.893392892893u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2271.802553053053u,0 2271.8035530530533u,1.5 2272.780093093093u,1.5 2272.781093093093u,0 2274.735173173173u,0 2274.736173173173u,1.5 2275.712713213213u,1.5 2275.7137132132134u,0 2276.690253253253u,0 2276.6912532532533u,1.5 2281.577953453453u,1.5 2281.5789534534533u,0 2285.488113613613u,0 2285.4891136136134u,1.5 2286.4656536536536u,1.5 2286.466653653654u,0 2287.4431936936935u,0 2287.4441936936937u,1.5 2288.420733733734u,1.5 2288.421733733734u,0 2289.3982737737733u,0 2289.3992737737735u,1.5 2291.3533538538536u,1.5 2291.354353853854u,0 2292.330893893894u,0 2292.331893893894u,1.5 2294.285973973974u,1.5 2294.286973973974u,0 2295.2635140140137u,0 2295.264514014014u,1.5 2296.241054054054u,1.5 2296.2420540540543u,0 2297.218594094094u,0 2297.219594094094u,1.5 2298.1961341341344u,1.5 2298.1971341341346u,0 2299.173674174174u,0 2299.174674174174u,1.5 2304.0613743743743u,1.5 2304.0623743743745u,0 2307.9715345345344u,0 2307.9725345345346u,1.5 2308.9490745745743u,1.5 2308.9500745745745u,0 2309.926614614614u,0 2309.9276146146144u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2317.746934934935u,0 2317.747934934935u,1.5 2319.7020150150147u,1.5 2319.703015015015u,0 2320.679555055055u,0 2320.6805550550553u,1.5 2326.5447952952954u,1.5 2326.5457952952956u,0 2329.477415415415u,0 2329.4784154154154u,1.5 2330.454955455455u,1.5 2330.4559554554553u,0 2331.4324954954955u,0 2331.4334954954957u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2343.1629759759758u,0 2343.163975975976u,1.5 2344.1405160160157u,1.5 2344.141516016016u,0 2346.095596096096u,0 2346.096596096096u,1.5 2347.0731361361363u,1.5 2347.0741361361365u,0 2349.028216216216u,0 2349.0292162162164u,1.5 2350.9832962962964u,1.5 2350.9842962962966u,0 2353.915916416416u,0 2353.9169164164164u,1.5 2355.8709964964964u,1.5 2355.8719964964966u,0 2356.8485365365364u,0 2356.8495365365366u,1.5 2357.8260765765763u,1.5 2357.8270765765765u,0 2359.7811566566565u,0 2359.7821566566568u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2361.736236736737u,0 2361.737236736737u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2365.646396896897u,1.5 2365.647396896897u,0 2368.5790170170167u,0 2368.580017017017u,1.5 2369.556557057057u,1.5 2369.5575570570572u,0 2370.534097097097u,0 2370.535097097097u,1.5 2371.5116371371373u,1.5 2371.5126371371375u,0 2372.4891771771768u,0 2372.490177177177u,1.5 2378.354417417417u,1.5 2378.3554174174174u,0 2379.331957457457u,0 2379.3329574574573u,1.5 2380.3094974974974u,1.5 2380.3104974974976u,0 2386.174737737738u,0 2386.175737737738u,1.5 2387.1522777777777u,1.5 2387.153277777778u,0 2390.084897897898u,0 2390.085897897898u,1.5 2392.039977977978u,1.5 2392.0409779779784u,0 2393.995058058058u,0 2393.996058058058u,1.5 2394.972598098098u,1.5 2394.973598098098u,0 2395.9501381381383u,0 2395.9511381381385u,1.5 2397.905218218218u,1.5 2397.9062182182183u,0 2398.882758258258u,0 2398.8837582582582u,1.5 2400.8378383383383u,1.5 2400.8388383383385u,0 2402.792918418418u,0 2402.7939184184183u,1.5 2403.7704584584585u,1.5 2403.7714584584587u,0 2404.7479984984984u,0 2404.7489984984986u,1.5 2406.7030785785787u,1.5 2406.704078578579u,0 2407.680618618618u,0 2407.6816186186184u,1.5 2408.6581586586585u,1.5 2408.6591586586587u,0 2409.6356986986984u,0 2409.6366986986986u,1.5 2413.5458588588585u,1.5 2413.5468588588587u,0 2419.411099099099u,0 2419.412099099099u,1.5 2420.3886391391393u,1.5 2420.3896391391395u,0 2423.321259259259u,0 2423.322259259259u,1.5 2426.2538793793797u,1.5 2426.25487937938u,0 2427.231419419419u,0 2427.2324194194193u,1.5 2430.1640395395393u,1.5 2430.1650395395395u,0 2432.119119619619u,0 2432.1201196196193u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.0068198198196u,0 2437.00781981982u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2446.78222022022u,0 2446.7832202202203u,1.5 2447.75976026026u,1.5 2447.76076026026u,0 2449.7148403403403u,0 2449.7158403403405u,1.5 2451.66992042042u,1.5 2451.6709204204203u,0 2452.6474604604605u,0 2452.6484604604607u,1.5 2453.6250005005004u,1.5 2453.6260005005006u,0 2454.6025405405403u,0 2454.6035405405405u,1.5 2463.400400900901u,1.5 2463.401400900901u,0 2465.355480980981u,0 2465.3564809809814u,1.5 2466.3330210210206u,1.5 2466.334021021021u,0 2467.310561061061u,0 2467.311561061061u,1.5 2469.2656411411413u,1.5 2469.2666411411415u,0 2470.243181181181u,0 2470.2441811811814u,1.5 2472.198261261261u,1.5 2472.199261261261u,0 2473.1758013013014u,0 2473.1768013013016u,1.5 2475.1308813813816u,1.5 2475.131881381382u,0 2476.108421421421u,0 2476.1094214214213u,1.5 2477.0859614614615u,1.5 2477.0869614614617u,0 2479.0410415415413u,0 2479.0420415415415u,1.5 2480.996121621621u,1.5 2480.9971216216213u,0 2484.9062817817817u,0 2484.907281781782u,1.5 2485.8838218218216u,1.5 2485.884821821822u,0 2487.838901901902u,0 2487.839901901902u,1.5 2489.793981981982u,1.5 2489.7949819819823u,0 2494.681682182182u,0 2494.6826821821824u,1.5 2495.659222222222u,1.5 2495.6602222222223u,0 2502.5020025025024u,0 2502.5030025025026u,1.5 2505.434622622622u,1.5 2505.4356226226223u,0 2507.3897027027024u,0 2507.3907027027026u,1.5 2508.3672427427427u,1.5 2508.368242742743u,0 2511.2998628628625u,0 2511.3008628628627u,1.5 2512.277402902903u,1.5 2512.278402902903u,0 2513.2549429429428u,0 2513.255942942943u,1.5 2516.187563063063u,1.5 2516.188563063063u,0 2522.0528033033033u,0 2522.0538033033035u,1.5 2523.0303433433432u,1.5 2523.0313433433435u,0 2524.0078833833836u,0 2524.008883383384u,1.5 2524.985423423423u,1.5 2524.9864234234233u,0 2526.9405035035034u,0 2526.9415035035036u,1.5 2527.9180435435437u,1.5 2527.919043543544u,0 2528.8955835835836u,0 2528.896583583584u,1.5 2530.8506636636635u,1.5 2530.8516636636637u,0 2531.8282037037034u,0 2531.8292037037036u,1.5 2532.8057437437437u,1.5 2532.806743743744u,0 2533.7832837837836u,0 2533.784283783784u,1.5 2535.7383638638635u,1.5 2535.7393638638637u,0 2536.715903903904u,0 2536.716903903904u,1.5 2538.670983983984u,1.5 2538.6719839839843u,0 2539.6485240240236u,0 2539.649524024024u,1.5 2540.626064064064u,1.5 2540.627064064064u,0 2542.581144144144u,0 2542.5821441441444u,1.5 2545.513764264264u,1.5 2545.514764264264u,0 2546.4913043043043u,0 2546.4923043043045u,1.5 2549.423924424424u,1.5 2549.4249244244243u,0 2550.4014644644644u,0 2550.4024644644646u,1.5 2552.3565445445447u,1.5 2552.357544544545u,0 2556.2667047047044u,0 2556.2677047047046u,1.5 2557.2442447447447u,1.5 2557.245244744745u,0 2559.1993248248245u,0 2559.2003248248247u,1.5 2560.1768648648645u,1.5 2560.1778648648647u,0 2563.109484984985u,0 2563.1104849849853u,1.5 2564.0870250250246u,1.5 2564.0880250250248u,0 2566.042105105105u,0 2566.043105105105u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2572.8848853853856u,0 2572.885885385386u,1.5 2574.8399654654654u,1.5 2574.8409654654656u,0 2575.8175055055053u,0 2575.8185055055055u,1.5 2577.7725855855856u,1.5 2577.773585585586u,0 2579.7276656656654u,0 2579.7286656656656u,1.5 2582.6602857857856u,1.5 2582.661285785786u,0 2583.6378258258255u,0 2583.6388258258257u,1.5 2584.6153658658654u,1.5 2584.6163658658656u,0 2588.5255260260255u,0 2588.5265260260257u,1.5 2590.480606106106u,1.5 2590.481606106106u,0 2593.413226226226u,0 2593.414226226226u,1.5 2594.390766266266u,1.5 2594.391766266266u,0 2595.3683063063063u,0 2595.3693063063065u,1.5 2597.3233863863866u,1.5 2597.324386386387u,0 2598.300926426426u,0 2598.3019264264262u,1.5 2599.2784664664664u,1.5 2599.2794664664666u,0 2600.2560065065063u,0 2600.2570065065065u,1.5 2602.2110865865866u,1.5 2602.212086586587u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2607.0987867867866u,0 2607.099786786787u,1.5 2613.941567067067u,1.5 2613.942567067067u,0 2617.851727227227u,0 2617.852727227227u,1.5 2618.829267267267u,1.5 2618.830267267267u,0 2620.784347347347u,0 2620.7853473473474u,1.5 2623.7169674674674u,1.5 2623.7179674674676u,0 2627.6271276276275u,0 2627.6281276276277u,1.5 2630.5597477477477u,1.5 2630.560747747748u,0 2636.424987987988u,0 2636.4259879879883u,1.5 2638.380068068068u,1.5 2638.381068068068u,0 2639.357608108108u,0 2639.358608108108u,1.5 2643.267768268268u,1.5 2643.268768268268u,0 2648.1554684684684u,0 2648.1564684684686u,1.5 2649.1330085085083u,1.5 2649.1340085085085u,0 2650.1105485485486u,0 2650.111548548549u,1.5 2652.065628628629u,1.5 2652.066628628629u,0 2653.0431686686684u,0 2653.0441686686686u,1.5 2654.0207087087088u,1.5 2654.021708708709u,0 2654.9982487487487u,0 2654.999248748749u,1.5 2655.9757887887886u,1.5 2655.976788788789u,0 2656.953328828829u,0 2656.954328828829u,1.5 2657.9308688688684u,1.5 2657.9318688688686u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2668.6838093093093u,1.5 2668.6848093093095u,0 2673.5715095095093u,0 2673.5725095095095u,1.5 2674.5490495495496u,1.5 2674.55004954955u,0 2676.50412962963u,0 2676.50512962963u,1.5 2677.4816696696694u,1.5 2677.4826696696696u,0 2678.4592097097097u,0 2678.46020970971u,1.5 2679.4367497497497u,1.5 2679.43774974975u,0 2680.4142897897896u,0 2680.4152897897898u,1.5 2681.39182982983u,1.5 2681.39282982983u,0 2686.27953003003u,0 2686.28053003003u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2689.21215015015u,1.5 2689.2131501501503u,0 2690.18969019019u,0 2690.1906901901903u,1.5 2692.14477027027u,1.5 2692.14577027027u,0 2694.09985035035u,0 2694.1008503503504u,1.5 2695.0773903903905u,1.5 2695.0783903903907u,0 2698.0100105105103u,0 2698.0110105105105u,1.5 2698.9875505505506u,1.5 2698.988550550551u,0 2699.9650905905905u,0 2699.9660905905907u,1.5 2700.942630630631u,1.5 2700.943630630631u,0 2701.9201706706704u,0 2701.9211706706706u,1.5 2702.8977107107107u,1.5 2702.898710710711u,0 2704.8527907907906u,0 2704.8537907907908u,1.5 2705.830330830831u,1.5 2705.831330830831u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2708.7629509509507u,1.5 2708.763950950951u,0 2709.740490990991u,0 2709.741490990991u,1.5 2710.718031031031u,1.5 2710.719031031031u,0 2711.695571071071u,0 2711.696571071071u,1.5 2712.6731111111108u,1.5 2712.674111111111u,0 2713.650651151151u,0 2713.6516511511513u,1.5 2714.628191191191u,1.5 2714.6291911911912u,0 2716.583271271271u,0 2716.584271271271u,1.5 2718.538351351351u,1.5 2718.5393513513513u,0 2719.5158913913915u,0 2719.5168913913917u,1.5 2721.4709714714713u,1.5 2721.4719714714715u,0 2723.4260515515516u,0 2723.427051551552u,1.5 2724.4035915915915u,1.5 2724.4045915915917u,0 2725.381131631632u,0 2725.382131631632u,1.5 2727.3362117117117u,1.5 2727.337211711712u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2732.2239119119117u,0 2732.224911911912u,1.5 2737.1116121121117u,1.5 2737.112612112112u,0 2739.066692192192u,0 2739.067692192192u,1.5 2740.0442322322324u,1.5 2740.0452322322326u,0 2741.021772272272u,0 2741.022772272272u,1.5 2745.9094724724723u,1.5 2745.9104724724725u,0 2749.819632632633u,0 2749.820632632633u,1.5 2755.6848728728723u,1.5 2755.6858728728726u,0 2757.6399529529526u,0 2757.640952952953u,1.5 2759.595033033033u,1.5 2759.596033033033u,0 2760.572573073073u,0 2760.573573073073u,1.5 2763.505193193193u,1.5 2763.506193193193u,0 2765.460273273273u,0 2765.461273273273u,1.5 2766.437813313313u,1.5 2766.4388133133134u,0 2768.3928933933935u,0 2768.3938933933937u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2775.2356736736733u,1.5 2775.2366736736735u,0 2777.1907537537536u,0 2777.191753753754u,1.5 2778.168293793794u,1.5 2778.169293793794u,0 2782.0784539539536u,0 2782.079453953954u,1.5 2785.9886141141137u,1.5 2785.989614114114u,0 2786.966154154154u,0 2786.9671541541543u,1.5 2787.943694194194u,1.5 2787.944694194194u,0 2790.876314314314u,0 2790.8773143143144u,1.5 2791.853854354354u,1.5 2791.8548543543543u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2793.8089344344344u,1.5 2793.8099344344346u,0 2794.7864744744743u,0 2794.7874744744745u,1.5 2795.764014514514u,1.5 2795.7650145145144u,0 2796.7415545545546u,0 2796.7425545545548u,1.5 2797.7190945945945u,1.5 2797.7200945945947u,0 2804.561874874875u,0 2804.562874874875u,1.5 2807.494494994995u,1.5 2807.495494994995u,0 2814.337275275275u,0 2814.338275275275u,1.5 2822.1575955955955u,1.5 2822.1585955955957u,0 2828.022835835836u,0 2828.023835835836u,1.5 2830.9554559559556u,1.5 2830.956455955956u,0 2831.932995995996u,0 2831.933995995996u,1.5 2832.910536036036u,1.5 2832.911536036036u,0 2833.888076076076u,0 2833.889076076076u,1.5 2834.8656161161157u,1.5 2834.866616116116u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2841.7083963963964u,1.5 2841.7093963963966u,0 2842.6859364364364u,0 2842.6869364364366u,1.5 2844.641016516516u,1.5 2844.6420165165164u,0 2845.6185565565565u,0 2845.6195565565567u,1.5 2849.5287167167166u,1.5 2849.529716716717u,0 2850.5062567567566u,0 2850.5072567567568u,1.5 2851.483796796797u,1.5 2851.484796796797u,0 2852.461336836837u,0 2852.462336836837u,1.5 2856.371496996997u,1.5 2856.372496996997u,0 2857.349037037037u,0 2857.350037037037u,1.5 2858.3265770770768u,1.5 2858.327577077077u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2864.191817317317u,0 2864.1928173173173u,1.5 2868.1019774774772u,1.5 2868.1029774774775u,0 2869.079517517517u,0 2869.0805175175174u,1.5 2870.0570575575575u,1.5 2870.0580575575577u,0 2871.0345975975974u,0 2871.0355975975976u,1.5 2872.012137637638u,1.5 2872.013137637638u,0 2876.899837837838u,0 2876.900837837838u,1.5 2877.877377877878u,1.5 2877.8783778778784u,0 2878.8549179179176u,0 2878.855917917918u,1.5 2880.809997997998u,1.5 2880.810997997998u,0 2883.7426181181177u,0 2883.743618118118u,1.5 2885.697698198198u,1.5 2885.698698198198u,0 2886.6752382382383u,0 2886.6762382382385u,1.5 2887.652778278278u,1.5 2887.6537782782784u,0 2888.630318318318u,0 2888.6313183183183u,1.5 2891.5629384384383u,1.5 2891.5639384384385u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2897.4281786786787u,1.5 2897.429178678679u,0 2898.4057187187186u,0 2898.406718718719u,1.5 2901.338338838839u,1.5 2901.339338838839u,0 2906.226039039039u,0 2906.227039039039u,1.5 2908.1811191191186u,1.5 2908.182119119119u,0 2911.1137392392393u,0 2911.1147392392395u,1.5 2912.091279279279u,1.5 2912.0922792792794u,0 2913.068819319319u,0 2913.0698193193193u,1.5 2917.956519519519u,1.5 2917.9575195195193u,0 2920.88913963964u,0 2920.89013963964u,1.5 2921.8666796796797u,1.5 2921.86767967968u,0 2922.8442197197196u,0 2922.84521971972u,1.5 2923.8217597597595u,1.5 2923.8227597597597u,0 2925.77683983984u,0 2925.77783983984u,1.5 2926.75437987988u,1.5 2926.7553798798804u,0 2927.7319199199196u,0 2927.73291991992u,1.5 2929.687u,1.5 2929.688u,0 2931.64208008008u,0 2931.6430800800804u,1.5 2932.6196201201196u,1.5 2932.62062012012u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2936.52978028028u,1.5 2936.5307802802804u,0 2937.50732032032u,0 2937.5083203203203u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2942.39502052052u,1.5 2942.3960205205203u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 2948.2602607607605u,1.5 2948.2612607607607u,0 2949.237800800801u,0 2949.238800800801u,1.5 2950.215340840841u,1.5 2950.216340840841u,0 2952.1704209209206u,0 2952.171420920921u,1.5 2953.147960960961u,1.5 2953.148960960961u,0 2955.103041041041u,0 2955.104041041041u,1.5 2957.0581211211206u,1.5 2957.059121121121u,0 2958.035661161161u,0 2958.036661161161u,1.5 2959.013201201201u,1.5 2959.014201201201u,0 2960.968281281281u,0 2960.9692812812814u,1.5 2966.833521521521u,1.5 2966.8345215215213u,0 2967.8110615615615u,0 2967.8120615615617u,1.5 2968.7886016016014u,1.5 2968.7896016016016u,0 2969.7661416416418u,0 2969.767141641642u,1.5 2970.7436816816817u,1.5 2970.744681681682u,0 2972.6987617617615u,0 2972.6997617617617u,1.5 2974.6538418418418u,1.5 2974.654841841842u,0 2975.631381881882u,0 2975.6323818818823u,1.5 2980.519082082082u,1.5 2980.5200820820824u,0 2981.4966221221216u,0 2981.497622122122u,1.5 2983.451702202202u,1.5 2983.452702202202u,0 2984.4292422422423u,0 2984.4302422422425u,1.5 2986.384322322322u,1.5 2986.3853223223223u,0 2988.3394024024024u,0 2988.3404024024026u,1.5 2989.3169424424423u,1.5 2989.3179424424425u,0 2990.2944824824826u,0 2990.295482482483u,1.5 2993.2271026026024u,1.5 2993.2281026026026u,0 2994.2046426426427u,0 2994.205642642643u,1.5 2997.1372627627625u,1.5 2997.1382627627627u,0 2998.114802802803u,0 2998.115802802803u,1.5 2999.0923428428428u,1.5 2999.093342842843u,0 3000.069882882883u,0 3000.0708828828833u,1.5 3003.980043043043u,1.5 3003.9810430430434u,0 3004.957583083083u,0 3004.9585830830833u,1.5 3010.822823323323u,1.5 3010.8238233233233u,0 3011.800363363363u,0 3011.801363363363u,1.5 3014.7329834834836u,1.5 3014.733983483484u,0 3015.710523523523u,0 3015.7115235235233u,1.5 3017.6656036036034u,1.5 3017.6666036036036u,0 3018.6431436436437u,0 3018.644143643644u,1.5 3022.553303803804u,1.5 3022.554303803804u,0 3023.5308438438437u,0 3023.531843843844u,1.5 3026.463463963964u,1.5 3026.464463963964u,0 3027.441004004004u,0 3027.442004004004u,1.5 3028.418544044044u,1.5 3028.4195440440444u,0 3029.396084084084u,0 3029.3970840840843u,1.5 3030.373624124124u,1.5 3030.3746241241242u,0 3032.328704204204u,0 3032.329704204204u,1.5 3033.306244244244u,1.5 3033.3072442442444u,0 3036.238864364364u,0 3036.239864364364u,1.5 3037.2164044044043u,1.5 3037.2174044044045u,0 3039.1714844844846u,0 3039.172484484485u,1.5 3040.149024524524u,1.5 3040.1500245245243u,0 3043.0816446446447u,0 3043.082644644645u,1.5 3044.0591846846846u,1.5 3044.060184684685u,0 3046.0142647647644u,0 3046.0152647647647u,1.5 3046.991804804805u,1.5 3046.992804804805u,0 3048.946884884885u,0 3048.9478848848853u,1.5 3050.901964964965u,1.5 3050.902964964965u,0 3051.879505005005u,0 3051.880505005005u,1.5 3059.699825325325u,1.5 3059.7008253253252u,0 3061.6549054054053u,0 3061.6559054054055u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3064.587525525525u,0 3064.5885255255253u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3069.4752257257255u,0 3069.4762257257257u,1.5 3070.4527657657654u,1.5 3070.4537657657656u,0 3073.385385885886u,0 3073.3863858858863u,1.5 3076.318006006006u,1.5 3076.319006006006u,0 3077.295546046046u,0 3077.2965460460464u,1.5 3081.205706206206u,1.5 3081.206706206206u,0 3082.183246246246u,0 3082.1842462462464u,1.5 3085.115866366366u,1.5 3085.116866366366u,0 3086.0934064064063u,0 3086.0944064064065u,1.5 3089.026026526526u,1.5 3089.0270265265262u,0 3093.9137267267265u,0 3093.9147267267267u,1.5 3094.8912667667664u,1.5 3094.8922667667666u,0 3096.8463468468467u,0 3096.847346846847u,1.5 3097.823886886887u,1.5 3097.8248868868873u,0 3100.756507007007u,0 3100.757507007007u,1.5 3102.711587087087u,1.5 3102.7125870870873u,0 3103.689127127127u,0 3103.690127127127u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3108.576827327327u,0 3108.577827327327u,1.5 3109.554367367367u,1.5 3109.555367367367u,0 3112.4869874874876u,0 3112.4879874874878u,1.5 3113.464527527527u,1.5 3113.4655275275272u,0 3114.4420675675674u,0 3114.4430675675676u,1.5 3119.3297677677674u,1.5 3119.3307677677676u,0 3121.2848478478477u,0 3121.285847847848u,1.5 3122.262387887888u,1.5 3122.2633878878883u,0 3128.127628128128u,0 3128.128628128128u,1.5 3129.105168168168u,1.5 3129.106168168168u,0 3130.0827082082083u,0 3130.0837082082085u,1.5 3132.037788288288u,1.5 3132.0387882882883u,0 3133.992868368368u,0 3133.993868368368u,1.5 3134.9704084084083u,1.5 3134.9714084084085u,0 3136.9254884884886u,0 3136.9264884884888u,1.5 3137.9030285285285u,1.5 3137.9040285285287u,0 3139.8581086086083u,0 3139.8591086086085u,1.5 3140.8356486486487u,1.5 3140.836648648649u,0 3141.8131886886886u,0 3141.814188688689u,1.5 3142.790728728729u,1.5 3142.791728728729u,0 3143.7682687687684u,0 3143.7692687687686u,1.5 3144.7458088088088u,1.5 3144.746808808809u,0 3146.700888888889u,0 3146.7018888888892u,1.5 3147.678428928929u,1.5 3147.679428928929u,0 3148.655968968969u,0 3148.656968968969u,1.5 3149.633509009009u,1.5 3149.634509009009u,0 3151.588589089089u,0 3151.5895890890893u,1.5 3153.543669169169u,1.5 3153.544669169169u,0 3154.5212092092092u,0 3154.5222092092094u,1.5 3155.498749249249u,1.5 3155.4997492492494u,0 3157.4538293293294u,0 3157.4548293293296u,1.5 3160.386449449449u,1.5 3160.3874494494494u,0 3162.3415295295295u,0 3162.3425295295297u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3164.2966096096093u,0 3164.2976096096095u,1.5 3166.2516896896896u,1.5 3166.2526896896898u,0 3168.2067697697694u,0 3168.2077697697696u,1.5 3169.1843098098097u,1.5 3169.18530980981u,0 3170.1618498498497u,0 3170.16284984985u,1.5 3174.0720100100098u,1.5 3174.07301001001u,0 3175.04955005005u,0 3175.0505500500503u,1.5 3176.02709009009u,1.5 3176.0280900900902u,0 3177.98217017017u,0 3177.98317017017u,1.5 3178.9597102102102u,1.5 3178.9607102102104u,0 3179.93725025025u,0 3179.9382502502503u,1.5 3180.91479029029u,1.5 3180.9157902902903u,0 3181.8923303303304u,0 3181.8933303303306u,1.5 3183.8474104104102u,1.5 3183.8484104104105u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3187.7575705705704u,1.5 3187.7585705705706u,0 3190.6901906906905u,0 3190.6911906906907u,1.5 3191.667730730731u,1.5 3191.668730730731u,0 3192.6452707707704u,0 3192.6462707707706u,1.5 3195.577890890891u,1.5 3195.578890890891u,0 3196.555430930931u,0 3196.556430930931u,1.5 3197.532970970971u,1.5 3197.533970970971u,0 3203.398211211211u,0 3203.3992112112114u,1.5 3204.375751251251u,1.5 3204.3767512512513u,0 3205.353291291291u,0 3205.3542912912912u,1.5 3209.263451451451u,1.5 3209.2644514514514u,0 3213.1736116116112u,0 3213.1746116116115u,1.5 3214.1511516516516u,1.5 3214.152151651652u,0 3217.0837717717714u,0 3217.0847717717716u,1.5 3218.0613118118117u,1.5 3218.062311811812u,0 3219.0388518518516u,0 3219.039851851852u,1.5 3220.016391891892u,1.5 3220.017391891892u,0 3223.926552052052u,0 3223.9275520520523u,1.5 3224.904092092092u,1.5 3224.905092092092u,0 3225.8816321321324u,0 3225.8826321321326u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3234.6794924924925u,0 3234.6804924924927u,1.5 3238.5896526526526u,1.5 3238.590652652653u,0 3240.544732732733u,0 3240.545732732733u,1.5 3241.5222727727723u,1.5 3241.5232727727725u,0 3244.454892892893u,0 3244.455892892893u,1.5 3246.409972972973u,1.5 3246.410972972973u,0 3247.3875130130127u,0 3247.388513013013u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3254.2302932932935u,0 3254.2312932932937u,1.5 3261.0730735735733u,1.5 3261.0740735735735u,0 3262.050613613613u,0 3262.0516136136134u,1.5 3263.0281536536536u,1.5 3263.029153653654u,0 3264.983233733734u,0 3264.984233733734u,1.5 3266.9383138138137u,1.5 3266.939313813814u,0 3267.9158538538536u,0 3267.916853853854u,1.5 3269.870933933934u,1.5 3269.871933933934u,0 3270.848473973974u,0 3270.849473973974u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3273.781094094094u,1.5 3273.782094094094u,0 3276.713714214214u,0 3276.7147142142144u,1.5 3280.6238743743743u,1.5 3280.6248743743745u,0 3281.601414414414u,0 3281.6024144144144u,1.5 3283.5564944944945u,1.5 3283.5574944944947u,0 3287.4666546546546u,0 3287.467654654655u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3297.242055055055u,0 3297.2430550550553u,1.5 3298.219595095095u,1.5 3298.220595095095u,0 3299.1971351351353u,0 3299.1981351351355u,1.5 3300.174675175175u,1.5 3300.175675175175u,0 3306.039915415415u,0 3306.0409154154154u,1.5 3307.017455455455u,1.5 3307.0184554554553u,0 3307.9949954954955u,0 3307.9959954954957u,1.5 3309.9500755755753u,1.5 3309.9510755755755u,0 3310.927615615615u,0 3310.9286156156154u,1.5 3312.8826956956955u,1.5 3312.8836956956957u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3315.8153158158157u,1.5 3315.816315815816u,0 3317.770395895896u,0 3317.771395895896u,1.5 3318.747935935936u,1.5 3318.748935935936u,0 3319.7254759759758u,0 3319.726475975976u,1.5 3323.6356361361363u,1.5 3323.6366361361365u,0 3324.613176176176u,0 3324.614176176176u,1.5 3325.590716216216u,1.5 3325.5917162162164u,0 3326.568256256256u,0 3326.5692562562563u,1.5 3330.478416416416u,1.5 3330.4794164164164u,0 3331.455956456456u,0 3331.4569564564563u,1.5 3332.4334964964964u,1.5 3332.4344964964966u,0 3333.4110365365364u,0 3333.4120365365366u,1.5 3335.366116616616u,1.5 3335.3671166166164u,0 3337.3211966966965u,0 3337.3221966966967u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3342.208896896897u,0 3342.209896896897u,1.5 3343.186436936937u,1.5 3343.187436936937u,0 3346.119057057057u,0 3346.1200570570572u,1.5 3350.029217217217u,1.5 3350.0302172172173u,0 3351.006757257257u,0 3351.0077572572573u,1.5 3351.9842972972974u,1.5 3351.9852972972976u,0 3355.894457457457u,0 3355.8954574574573u,1.5 3356.8719974974974u,1.5 3356.8729974974976u,0 3357.8495375375373u,0 3357.8505375375375u,1.5 3360.7821576576575u,1.5 3360.7831576576577u,0 3363.7147777777773u,0 3363.7157777777775u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3369.5800180180177u,0 3369.581018018018u,1.5 3371.535098098098u,1.5 3371.536098098098u,0 3372.5126381381383u,0 3372.5136381381385u,1.5 3373.4901781781778u,1.5 3373.491178178178u,0 3374.467718218218u,0 3374.4687182182183u,1.5 3379.355418418418u,1.5 3379.3564184184183u,0 3382.2880385385383u,0 3382.2890385385385u,1.5 3383.2655785785787u,1.5 3383.266578578579u,0 3386.1981986986984u,0 3386.1991986986986u,1.5 3387.175738738739u,1.5 3387.176738738739u,0 3390.1083588588585u,0 3390.1093588588587u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.0185190190186u,0 3394.019519019019u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3398.906219219219u,0 3398.9072192192193u,1.5 3399.883759259259u,1.5 3399.884759259259u,0 3400.8612992992994u,0 3400.8622992992996u,1.5 3401.8388393393393u,1.5 3401.8398393393395u,0 3403.793919419419u,0 3403.7949194194193u,1.5 3407.7040795795797u,1.5 3407.70507957958u,0 3409.6591596596595u,0 3409.6601596596597u,1.5 3410.6366996996994u,1.5 3410.6376996996996u,0 3411.61423973974u,0 3411.61523973974u,1.5 3412.5917797797797u,1.5 3412.59277977978u,0 3414.5468598598595u,0 3414.5478598598597u,1.5 3415.5243998999u,1.5 3415.5253998999u,0 3420.4121001001u,0 3420.4131001001u,1.5 3421.3896401401403u,1.5 3421.3906401401405u,0 3422.36718018018u,0 3422.3681801801804u,1.5 3424.32226026026u,1.5 3424.32326026026u,0 3425.2998003003004u,0 3425.3008003003006u,1.5 3427.2548803803807u,1.5 3427.255880380381u,0 3428.23242042042u,0 3428.2334204204203u,1.5 3429.2099604604605u,1.5 3429.2109604604607u,0 3430.1875005005004u,0 3430.1885005005006u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3437.0302807807807u,1.5 3437.031280780781u,0 3438.0078208208206u,0 3438.008820820821u,1.5 3438.9853608608605u,1.5 3438.9863608608607u,0 3446.805681181181u,0 3446.8066811811814u,1.5 3447.783221221221u,1.5 3447.7842212212213u,0 3450.7158413413413u,0 3450.7168413413415u,1.5 3452.670921421421u,1.5 3452.6719214214213u,0 3453.6484614614615u,0 3453.6494614614617u,1.5 3454.6260015015014u,1.5 3454.6270015015016u,0 3456.5810815815817u,0 3456.582081581582u,1.5 3460.4912417417418u,1.5 3460.492241741742u,0 3461.4687817817817u,0 3461.469781781782u,1.5 3465.378941941942u,1.5 3465.379941941942u,0 3466.356481981982u,0 3466.3574819819823u,1.5 3467.3340220220216u,1.5 3467.335022022022u,0 3468.311562062062u,0 3468.312562062062u,1.5 3469.289102102102u,1.5 3469.290102102102u,0 3470.2666421421422u,0 3470.2676421421424u,1.5 3472.221722222222u,1.5 3472.2227222222223u,0 3473.199262262262u,0 3473.200262262262u,1.5 3474.1768023023023u,1.5 3474.1778023023026u,0 3475.1543423423423u,0 3475.1553423423425u,1.5 3476.1318823823826u,1.5 3476.132882382383u,0 3478.0869624624625u,0 3478.0879624624627u,1.5 3479.0645025025024u,1.5 3479.0655025025026u,0 3481.0195825825826u,0 3481.020582582583u,1.5 3481.997122622622u,1.5 3481.9981226226223u,0 3482.9746626626625u,0 3482.9756626626627u,1.5 3483.9522027027024u,1.5 3483.9532027027026u,0 3493.727603103103u,0 3493.728603103103u,1.5 3494.7051431431432u,1.5 3494.7061431431434u,0 3495.682683183183u,0 3495.6836831831833u,1.5 3496.660223223223u,1.5 3496.6612232232233u,0 3501.547923423423u,0 3501.5489234234233u,1.5 3503.5030035035034u,1.5 3503.5040035035036u,0 3521.098724224224u,0 3521.0997242242242u,1.5 3522.076264264264u,1.5 3522.077264264264u,0 3525.0088843843846u,0 3525.009884384385u,1.5 3526.9639644644644u,1.5 3526.9649644644646u,0 3527.9415045045043u,0 3527.9425045045045u,1.5 3529.8965845845846u,1.5 3529.897584584585u,0 3530.8741246246245u,0 3530.8751246246247u,1.5 3531.8516646646644u,1.5 3531.8526646646646u,0 3533.8067447447447u,0 3533.807744744745u,1.5 3535.7618248248245u,1.5 3535.7628248248247u,0 3536.7393648648645u,0 3536.7403648648647u,1.5 3537.716904904905u,1.5 3537.717904904905u,0 3539.671984984985u,0 3539.6729849849853u,1.5 3540.6495250250246u,1.5 3540.6505250250248u,0 3541.627065065065u,0 3541.628065065065u,1.5 3542.604605105105u,1.5 3542.605605105105u,0 3543.582145145145u,0 3543.5831451451454u,1.5 3546.514765265265u,1.5 3546.515765265265u,0 3547.4923053053053u,0 3547.4933053053055u,1.5 3548.469845345345u,1.5 3548.4708453453454u,0 3549.4473853853856u,0 3549.448385385386u,1.5 3551.4024654654654u,1.5 3551.4034654654656u,0 3553.3575455455457u,0 3553.358545545546u,1.5 3554.3350855855856u,1.5 3554.336085585586u,0 3555.3126256256255u,0 3555.3136256256257u,1.5 3556.2901656656654u,1.5 3556.2911656656656u,0 3561.1778658658654u,0 3561.1788658658656u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3564.110485985986u,0 3564.1114859859863u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.998186186186u,1.5 3568.9991861861863u,0 3570.953266266266u,0 3570.954266266266u,1.5 3574.863426426426u,1.5 3574.8644264264262u,0 3576.8185065065063u,0 3576.8195065065065u,1.5 3577.7960465465467u,1.5 3577.797046546547u,0 3578.7735865865866u,0 3578.774586586587u,1.5 3579.7511266266265u,1.5 3579.7521266266267u,0 3581.7062067067063u,0 3581.7072067067065u,1.5 3582.6837467467467u,1.5 3582.684746746747u,0 3583.6612867867866u,0 3583.662286786787u,1.5 3584.6388268268265u,1.5 3584.6398268268267u,0 3586.593906906907u,0 3586.594906906907u,1.5 3588.548986986987u,1.5 3588.5499869869873u,0 3589.5265270270265u,0 3589.5275270270267u,1.5 3597.346847347347u,1.5 3597.3478473473474u,0 3598.3243873873876u,0 3598.3253873873878u,1.5 3599.301927427427u,1.5 3599.302927427427u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3609.0773278278275u,0 3609.0783278278277u,1.5 3612.0099479479477u,1.5 3612.010947947948u,0 3612.987487987988u,0 3612.9884879879883u,1.5 3613.9650280280275u,1.5 3613.9660280280277u,0 3615.920108108108u,0 3615.921108108108u,1.5 3616.897648148148u,1.5 3616.8986481481484u,0 3617.875188188188u,0 3617.8761881881883u,1.5 3619.830268268268u,1.5 3619.831268268268u,0 3621.785348348348u,0 3621.7863483483484u,1.5 3622.7628883883885u,1.5 3622.7638883883888u,0 3623.740428428428u,0 3623.741428428428u,1.5 3624.7179684684684u,1.5 3624.7189684684686u,0 3625.6955085085083u,0 3625.6965085085085u,1.5 3627.6505885885886u,1.5 3627.6515885885888u,0 3628.6281286286285u,0 3628.6291286286287u,1.5 3630.5832087087088u,1.5 3630.584208708709u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3640.358609109109u,1.5 3640.359609109109u,0 3641.336149149149u,0 3641.3371491491494u,1.5 3643.2912292292294u,1.5 3643.2922292292296u,0 3650.1340095095093u,0 3650.1350095095095u,1.5 3651.1115495495496u,1.5 3651.11254954955u,0 3652.0890895895895u,0 3652.0900895895898u,1.5 3655.9992497497497u,1.5 3656.00024974975u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3666.75219019019u,1.5 3666.7531901901903u,0 3667.7297302302304u,0 3667.7307302302306u,1.5 3670.66235035035u,1.5 3670.6633503503504u,0 3675.5500505505506u,0 3675.551050550551u,1.5 3676.5275905905905u,1.5 3676.5285905905907u,0 3677.505130630631u,0 3677.506130630631u,1.5 3678.4826706706704u,1.5 3678.4836706706706u,0 3679.4602107107107u,0 3679.461210710711u,1.5 3682.392830830831u,1.5 3682.393830830831u,0 3685.3254509509507u,0 3685.326450950951u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3689.2356111111108u,1.5 3689.236611111111u,0 3690.213151151151u,0 3690.2141511511513u,1.5 3691.190691191191u,1.5 3691.1916911911912u,0 3693.145771271271u,0 3693.146771271271u,1.5 3694.123311311311u,1.5 3694.1243113113114u,0 3697.0559314314314u,0 3697.0569314314316u,1.5 3698.0334714714713u,1.5 3698.0344714714715u,0 3699.0110115115112u,0 3699.0120115115114u,1.5 3702.9211716716713u,1.5 3702.9221716716715u,0 3703.8987117117117u,0 3703.899711711712u,1.5 3705.8537917917915u,1.5 3705.8547917917917u,0 3707.8088718718714u,0 3707.8098718718716u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3713.6741121121117u,1.5 3713.675112112112u,0 3718.561812312312u,0 3718.5628123123124u,1.5 3719.539352352352u,1.5 3719.5403523523523u,0 3720.5168923923925u,0 3720.5178923923927u,1.5 3723.4495125125122u,1.5 3723.4505125125124u,0 3725.4045925925925u,0 3725.4055925925927u,1.5 3726.382132632633u,1.5 3726.383132632633u,0 3728.3372127127127u,0 3728.338212712713u,1.5 3729.3147527527526u,1.5 3729.315752752753u,0 3730.292292792793u,0 3730.293292792793u,1.5 3732.2473728728723u,1.5 3732.2483728728726u,0 3735.179992992993u,0 3735.180992992993u,1.5 3736.157533033033u,1.5 3736.158533033033u,0 3740.067693193193u,0 3740.068693193193u,1.5 3744.9553933933935u,1.5 3744.9563933933937u,0 3745.9329334334334u,0 3745.9339334334336u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3755.708333833834u,1.5 3755.709333833834u,0 3758.6409539539536u,0 3758.641953953954u,1.5 3759.618493993994u,1.5 3759.619493993994u,0 3760.596034034034u,0 3760.597034034034u,1.5 3762.5511141141137u,1.5 3762.552114114114u,0 3764.506194194194u,0 3764.507194194194u,1.5 3766.461274274274u,1.5 3766.462274274274u,0 3770.3714344344344u,0 3770.3724344344346u,1.5 3775.259134634635u,1.5 3775.260134634635u,0 3776.2366746746743u,0 3776.2376746746745u,1.5 3778.1917547547546u,1.5 3778.192754754755u,0 3780.146834834835u,0 3780.147834834835u,1.5 3786.012075075075u,1.5 3786.013075075075u,0 3786.9896151151147u,0 3786.990615115115u,1.5 3787.967155155155u,1.5 3787.9681551551553u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3795.7874754754753u,1.5 3795.7884754754755u,0 3796.765015515515u,0 3796.7660155155154u,1.5 3797.7425555555556u,1.5 3797.7435555555558u,0 3799.697635635636u,0 3799.698635635636u,1.5 3801.6527157157157u,1.5 3801.653715715716u,0 3804.585335835836u,0 3804.586335835836u,1.5 3809.473036036036u,1.5 3809.474036036036u,0 3815.338276276276u,0 3815.339276276276u,1.5 3820.2259764764763u,1.5 3820.2269764764765u,0 3821.203516516516u,0 3821.2045165165164u,1.5 3822.1810565565565u,1.5 3822.1820565565567u,0 3829.023836836837u,0 3829.024836836837u,1.5 3830.9789169169167u,1.5 3830.979916916917u,0 3831.9564569569566u,0 3831.957456956957u,1.5 3833.911537037037u,1.5 3833.912537037037u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3839.776777277277u,1.5 3839.777777277277u,0 3840.754317317317u,0 3840.7553173173173u,1.5 3844.6644774774772u,1.5 3844.6654774774775u,0 3846.6195575575575u,0 3846.6205575575577u,1.5 3847.5970975975974u,1.5 3847.5980975975976u,0 3851.5072577577575u,0 3851.5082577577577u,1.5 3854.4398778778777u,1.5 3854.440877877878u,0 3855.4174179179176u,0 3855.418417917918u,1.5 3856.394957957958u,1.5 3856.395957957958u,0 3857.372497997998u,0 3857.373497997998u,1.5 3858.350038038038u,1.5 3858.351038038038u,0 3862.260198198198u,0 3862.261198198198u,1.5 3864.2152782782778u,1.5 3864.216278278278u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3870.080518518518u,1.5 3870.0815185185184u,0 3872.0355985985984u,0 3872.0365985985986u,1.5 3873.9906786786783u,1.5 3873.9916786786785u,0 3877.900838838839u,0 3877.901838838839u,1.5 3878.878378878879u,1.5 3878.8793788788794u,0 3879.8559189189186u,0 3879.856918918919u,1.5 3886.698699199199u,1.5 3886.699699199199u,0 3887.6762392392393u,0 3887.6772392392395u,1.5 3890.608859359359u,1.5 3890.6098593593592u,0 3892.5639394394393u,0 3892.5649394394395u,1.5 3903.31687987988u,1.5 3903.3178798798804u,0 3904.2944199199196u,0 3904.29541991992u,1.5 3905.27195995996u,1.5 3905.27295995996u,0 3907.22704004004u,0 3907.22804004004u,1.5 3908.20458008008u,1.5 3908.2055800800804u,0 3909.1821201201196u,0 3909.18312012012u,1.5 3910.1596601601605u,1.5 3910.1606601601607u,0 3913.09228028028u,0 3913.0932802802804u,1.5 3920.9126006006004u,1.5 3920.9136006006006u,0 3923.8452207207206u,0 3923.846220720721u,1.5 3924.822760760761u,1.5 3924.823760760761u,0 3928.7329209209206u,0 3928.733920920921u,1.5 3930.688001001001u,1.5 3930.689001001001u,0 3931.665541041041u,0 3931.666541041041u,1.5 3932.643081081081u,1.5 3932.6440810810814u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3937.530781281281u,0 3937.5317812812814u,1.5 3943.396021521521u,1.5 3943.3970215215213u,0 3944.373561561562u,0 3944.374561561562u,1.5 3947.3061816816817u,1.5 3947.307181681682u,0 3949.261261761762u,0 3949.262261761762u,1.5 3951.2163418418413u,1.5 3951.2173418418415u,0 3953.1714219219216u,0 3953.172421921922u,1.5 3954.1489619619624u,1.5 3954.1499619619626u,0 3955.126502002002u,0 3955.127502002002u,1.5 3956.104042042042u,1.5 3956.105042042042u,0 3957.081582082082u,0 3957.0825820820824u,1.5 3959.0366621621624u,1.5 3959.0376621621626u,0 3960.991742242242u,0 3960.992742242242u,1.5 3961.969282282282u,1.5 3961.9702822822824u,0 3964.9019024024024u,0 3964.9029024024026u,1.5 3965.879442442442u,1.5 3965.880442442442u,0 3966.8569824824826u,0 3966.857982482483u,1.5 3969.7896026026024u,1.5 3969.7906026026026u,0 3970.7671426426423u,0 3970.7681426426425u,1.5 3971.7446826826827u,1.5 3971.745682682683u,0 3972.7222227227226u,0 3972.7232227227228u,1.5 3974.677302802803u,1.5 3974.678302802803u,0 3976.632382882883u,0 3976.6333828828833u,1.5 3977.6099229229226u,1.5 3977.610922922923u,0 3978.5874629629634u,0 3978.5884629629636u,1.5 3985.430243243243u,1.5 3985.431243243243u,0 3986.407783283283u,0 3986.4087832832834u,1.5 3990.317943443443u,1.5 3990.318943443443u,0 3992.273023523523u,0 3992.2740235235233u,1.5 3994.2281036036034u,1.5 3994.2291036036036u,0 3995.2056436436433u,0 3995.2066436436435u,1.5 3996.1831836836836u,1.5 3996.184183683684u,0 3997.1607237237235u,0 3997.1617237237238u,1.5 3998.138263763764u,1.5 3998.139263763764u,0 4000.0933438438433u,0 4000.0943438438435u,1.5 4003.0259639639644u,1.5 4003.0269639639646u,0 4004.003504004004u,0 4004.004504004004u,1.5 4004.9810440440438u,1.5 4004.982044044044u,0 4005.958584084084u,0 4005.9595840840843u,1.5 4010.846284284284u,1.5 4010.8472842842843u,0 4013.7789044044043u,0 4013.7799044044045u,1.5 4018.6666046046043u,1.5 4018.6676046046045u,0 4019.6441446446443u,0 4019.6451446446445u,1.5 4023.554304804805u,1.5 4023.555304804805u,0 4024.5318448448443u,0 4024.5328448448445u,1.5 4025.509384884885u,1.5 4025.5103848848853u,0 4026.4869249249246u,0 4026.4879249249248u,1.5 4027.4644649649654u,1.5 4027.4654649649656u,0 4028.442005005005u,0 4028.443005005005u,1.5 4029.4195450450447u,1.5 4029.420545045045u,0 4031.374625125125u,0 4031.375625125125u,1.5 4032.3521651651654u,1.5 4032.3531651651656u,0 4033.329705205205u,0 4033.330705205205u,1.5 4035.284785285285u,1.5 4035.2857852852853u,0 4038.2174054054053u,0 4038.2184054054055u,1.5 4039.194945445445u,1.5 4039.195945445445u,0 4042.127565565566u,0 4042.128565565566u,1.5 4043.1051056056053u,1.5 4043.1061056056055u,0 4045.0601856856856u,0 4045.061185685686u,1.5 4046.0377257257255u,1.5 4046.0387257257257u,0 4047.992805805806u,0 4047.993805805806u,1.5 4048.9703458458453u,1.5 4048.9713458458455u,0 4049.947885885886u,0 4049.9488858858863u,1.5 4050.9254259259255u,1.5 4050.9264259259257u,0 4051.9029659659664u,0 4051.9039659659666u,1.5 4054.835586086086u,1.5 4054.8365860860863u,0 4055.813126126126u,0 4055.814126126126u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4072.431306806807u,1.5 4072.432306806807u,0 4075.3639269269265u,0 4075.3649269269267u,1.5 4077.319007007007u,1.5 4077.320007007007u,0 4080.251627127127u,0 4080.252627127127u,1.5 4081.2291671671674u,1.5 4081.2301671671676u,0 4083.1842472472467u,0 4083.185247247247u,1.5 4087.0944074074073u,1.5 4087.0954074074075u,0 4089.0494874874876u,0 4089.0504874874878u,1.5 4090.027027527527u,1.5 4090.0280275275272u,0 4093.9371876876876u,0 4093.938187687688u,1.5 4094.9147277277275u,1.5 4094.9157277277277u,0 4095.892267767768u,0 4095.893267767768u,1.5 4096.869807807808u,1.5 4096.870807807808u,0 4097.847347847847u,0 4097.848347847847u,1.5 4103.7125880880885u,1.5 4103.713588088089u,0 4104.690128128128u,0 4104.691128128128u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4111.532908408408u,0 4111.533908408408u,1.5 4112.510448448448u,1.5 4112.511448448448u,0 4113.487988488489u,0 4113.488988488489u,1.5 4120.330768768769u,1.5 4120.3317687687695u,0 4121.308308808809u,0 4121.309308808809u,1.5 4122.285848848848u,1.5 4122.286848848848u,0 4124.240928928929u,0 4124.241928928929u,1.5 4125.218468968969u,1.5 4125.2194689689695u,0 4129.128629129129u,0 4129.129629129129u,1.5 4130.106169169169u,1.5 4130.1071691691695u,0 4132.061249249249u,0 4132.062249249249u,1.5 4136.948949449449u,1.5 4136.949949449449u,0 4138.904029529529u,0 4138.905029529529u,1.5 4139.881569569569u,1.5 4139.88256956957u,0 4142.81418968969u,0 4142.81518968969u,1.5 4148.67942992993u,1.5 4148.68042992993u,0 4149.65696996997u,0 4149.6579699699705u,1.5 4150.63451001001u,1.5 4150.63551001001u,0 4154.54467017017u,0 4154.5456701701705u,1.5 4156.49975025025u,1.5 4156.50075025025u,0 4157.4772902902905u,0 4157.478290290291u,1.5 4160.40991041041u,1.5 4160.41091041041u,0 4161.38745045045u,0 4161.38845045045u,1.5 4162.3649904904905u,1.5 4162.365990490491u,0 4164.32007057057u,0 4164.321070570571u,1.5 4165.297610610611u,1.5 4165.298610610611u,0 4166.27515065065u,0 4166.27615065065u,1.5 4167.2526906906905u,1.5 4167.253690690691u,0 4168.23023073073u,0 4168.23123073073u,1.5 4172.140390890891u,1.5 4172.141390890891u,0 4178.005631131131u,0 4178.006631131131u,1.5 4178.983171171171u,1.5 4178.9841711711715u,0 4180.938251251251u,0 4180.939251251251u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4188.758571571571u,1.5 4188.7595715715715u,0 4191.6911916916915u,0 4191.692191691692u,1.5 4192.668731731731u,1.5 4192.669731731731u,0 4194.623811811812u,0 4194.624811811812u,1.5 4197.556431931932u,1.5 4197.557431931932u,0 4198.533971971972u,0 4198.5349719719725u,1.5 4199.511512012012u,1.5 4199.512512012012u,0 4200.489052052051u,0 4200.490052052051u,1.5 4201.4665920920925u,1.5 4201.467592092093u,0 4202.444132132132u,0 4202.445132132132u,1.5 4206.3542922922925u,1.5 4206.355292292293u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4210.264452452452u,0 4210.265452452452u,1.5 4212.219532532532u,1.5 4212.220532532532u,0 4213.197072572572u,0 4213.1980725725725u,1.5 4214.174612612613u,1.5 4214.175612612613u,0 4215.152152652652u,0 4215.153152652652u,1.5 4217.107232732732u,1.5 4217.108232732732u,0 4218.084772772773u,0 4218.085772772773u,1.5 4219.062312812813u,1.5 4219.063312812813u,0 4224.927553053052u,0 4224.928553053052u,1.5 4228.837713213213u,1.5 4228.838713213213u,0 4230.7927932932935u,0 4230.793793293294u,1.5 4231.770333333333u,1.5 4231.771333333333u,0 4234.702953453453u,0 4234.703953453453u,1.5 4236.658033533533u,1.5 4236.659033533533u,0 4238.613113613614u,0 4238.614113613614u,1.5 4240.5681936936935u,1.5 4240.569193693694u,0 4242.523273773774u,0 4242.524273773774u,1.5 4246.433433933934u,1.5 4246.434433933934u,0 4247.410973973974u,0 4247.411973973974u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4255.2312942942945u,0 4255.232294294295u,1.5 4256.208834334334u,1.5 4256.209834334334u,0 4257.186374374374u,0 4257.1873743743745u,1.5 4261.096534534534u,1.5 4261.097534534534u,0 4263.051614614615u,0 4263.052614614615u,1.5 4264.029154654655u,1.5 4264.030154654655u,0 4265.984234734734u,0 4265.985234734734u,1.5 4266.961774774775u,1.5 4266.962774774775u,0 4267.939314814815u,0 4267.940314814815u,1.5 4271.849474974975u,1.5 4271.850474974975u,0 4275.759635135135u,0 4275.760635135135u,1.5 4277.714715215215u,1.5 4277.715715215215u,0 4278.692255255256u,0 4278.693255255256u,1.5 4279.669795295295u,1.5 4279.670795295296u,0 4280.647335335335u,0 4280.648335335335u,1.5 4281.624875375375u,1.5 4281.6258753753755u,0 4284.5574954954955u,0 4284.558495495496u,1.5 4285.535035535535u,1.5 4285.536035535535u,0 4287.490115615616u,0 4287.491115615616u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4299.220596096096u,0 4299.221596096097u,1.5 4301.175676176176u,1.5 4301.176676176176u,0 4302.153216216216u,0 4302.154216216216u,1.5 4303.130756256257u,1.5 4303.131756256257u,0 4308.995996496496u,0 4308.996996496497u,1.5 4309.973536536536u,1.5 4309.974536536536u,0 4310.951076576576u,0 4310.9520765765765u,1.5 4315.838776776777u,1.5 4315.839776776777u,0 4316.816316816817u,0 4316.817316816817u,1.5 4317.793856856857u,1.5 4317.794856856857u,0 4318.7713968968965u,0 4318.772396896897u,1.5 4319.748936936937u,1.5 4319.749936936937u,0 4320.726476976977u,0 4320.727476976977u,1.5 4321.704017017017u,1.5 4321.705017017017u,0 4322.681557057057u,0 4322.682557057057u,1.5 4325.614177177177u,1.5 4325.615177177177u,0 4326.591717217217u,0 4326.592717217217u,1.5 4327.569257257258u,1.5 4327.570257257258u,0 4328.546797297297u,0 4328.547797297298u,1.5 4329.524337337337u,1.5 4329.525337337337u,0 4330.501877377377u,0 4330.502877377377u,1.5 4333.434497497497u,1.5 4333.435497497498u,0 4335.389577577577u,0 4335.3905775775775u,1.5 4338.322197697697u,1.5 4338.323197697698u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4342.232357857858u,0 4342.233357857858u,1.5 4344.187437937938u,1.5 4344.188437937938u,0 4345.164977977978u,0 4345.165977977978u,1.5 4351.030218218218u,1.5 4351.031218218218u,0 4352.007758258259u,0 4352.008758258259u,1.5 4352.985298298298u,1.5 4352.986298298299u,0 4353.962838338338u,0 4353.963838338338u,1.5 4354.940378378378u,1.5 4354.941378378378u,0 4357.872998498498u,0 4357.873998498499u,1.5 4358.850538538538u,1.5 4358.851538538538u,0 4359.828078578578u,0 4359.829078578578u,1.5 4360.805618618619u,1.5 4360.806618618619u,0 4361.783158658659u,0 4361.784158658659u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4371.558559059059u,0 4371.559559059059u,1.5 4374.491179179179u,1.5 4374.492179179179u,0 4375.468719219219u,0 4375.469719219219u,1.5 4376.44625925926u,1.5 4376.44725925926u,0 4377.423799299299u,0 4377.4247992993u,1.5 4379.378879379379u,1.5 4379.379879379379u,0 4384.266579579579u,0 4384.267579579579u,1.5 4387.199199699699u,1.5 4387.2001996997u,0 4388.176739739739u,0 4388.177739739739u,1.5 4389.15427977978u,1.5 4389.15527977978u,0 4390.13181981982u,0 4390.13281981982u,1.5 4392.086899899899u,1.5 4392.0878998999u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.01952002002u,0 4395.02052002002u,1.5 4397.95214014014u,1.5 4397.95314014014u,0 4402.83984034034u,0 4402.84084034034u,1.5 4403.81738038038u,1.5 4403.81838038038u,0 4405.772460460461u,0 4405.773460460461u,1.5 4407.72754054054u,1.5 4407.72854054054u,0 4408.70508058058u,0 4408.70608058058u,1.5 4409.682620620621u,1.5 4409.683620620621u,0 4410.660160660661u,0 4410.661160660661u,1.5 4412.61524074074u,1.5 4412.61624074074u,0 4414.570320820821u,0 4414.571320820821u,1.5 4415.547860860861u,1.5 4415.548860860861u,0 4417.502940940941u,0 4417.503940940941u,1.5 4418.480480980981u,1.5 4418.481480980981u,0 4422.390641141141u,0 4422.391641141141u,1.5 4424.345721221221u,1.5 4424.346721221221u,0 4425.323261261262u,0 4425.324261261262u,1.5 4426.300801301301u,1.5 4426.301801301302u,0 4427.278341341341u,0 4427.279341341341u,1.5 4430.210961461462u,1.5 4430.211961461462u,0 4431.188501501501u,0 4431.189501501502u,1.5 4432.166041541541u,1.5 4432.167041541541u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4439.008821821822u,0 4439.009821821822u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4443.896522022022u,0 4443.897522022022u,1.5 4444.874062062062u,1.5 4444.875062062062u,0 4446.829142142142u,0 4446.830142142142u,1.5 4448.784222222222u,1.5 4448.785222222222u,0 4449.761762262263u,0 4449.762762262263u,1.5 4450.739302302302u,1.5 4450.740302302303u,0 4451.716842342342u,0 4451.717842342342u,1.5 4453.6719224224225u,1.5 4453.672922422423u,0 4454.649462462463u,0 4454.650462462463u,1.5 4456.604542542542u,1.5 4456.605542542542u,0 4460.514702702702u,0 4460.515702702703u,1.5 4467.357482982983u,1.5 4467.358482982983u,0 4468.335023023023u,0 4468.336023023023u,1.5 4469.312563063063u,1.5 4469.313563063063u,0 4471.267643143143u,0 4471.268643143143u,1.5 4472.245183183183u,1.5 4472.246183183183u,0 4473.222723223223u,0 4473.223723223223u,1.5 4474.200263263264u,1.5 4474.201263263264u,0 4475.177803303303u,0 4475.1788033033035u,1.5 4476.155343343343u,1.5 4476.156343343343u,0 4478.1104234234235u,0 4478.111423423424u,1.5 4479.087963463464u,1.5 4479.088963463464u,0 4482.9981236236235u,0 4482.999123623624u,1.5 4485.930743743743u,1.5 4485.931743743743u,0 4491.795983983984u,0 4491.796983983984u,1.5 4492.773524024024u,1.5 4492.774524024024u,0 4494.728604104104u,0 4494.7296041041045u,1.5 4496.683684184184u,1.5 4496.684684184184u,0 4503.526464464465u,0 4503.527464464465u,1.5 4504.504004504504u,1.5 4504.5050045045045u,0 4505.481544544544u,0 4505.482544544544u,1.5 4508.414164664665u,1.5 4508.415164664665u,0 4510.369244744744u,0 4510.370244744744u,1.5 4511.346784784785u,1.5 4511.347784784785u,0 4514.279404904904u,0 4514.280404904905u,1.5 4515.256944944945u,1.5 4515.257944944945u,0 4519.167105105105u,0 4519.1681051051055u,1.5 4520.144645145145u,1.5 4520.145645145145u,0 4522.099725225225u,0 4522.100725225225u,1.5 4523.077265265266u,1.5 4523.078265265266u,0 4525.032345345345u,0 4525.033345345345u,1.5 4526.9874254254255u,1.5 4526.988425425426u,0 4528.942505505505u,0 4528.9435055055055u,1.5 4529.920045545545u,1.5 4529.921045545545u,0 4531.8751256256255u,0 4531.876125625626u,1.5 4536.7628258258255u,1.5 4536.763825825826u,0 4537.740365865866u,0 4537.741365865866u,1.5 4539.695445945946u,1.5 4539.696445945946u,0 4540.672985985986u,0 4540.673985985986u,1.5 4541.650526026026u,1.5 4541.651526026026u,0 4544.583146146146u,0 4544.584146146146u,1.5 4545.560686186186u,1.5 4545.561686186186u,0 4546.538226226226u,0 4546.539226226226u,1.5 4548.493306306306u,1.5 4548.4943063063065u,0 4550.448386386386u,0 4550.449386386386u,1.5 4551.4259264264265u,1.5 4551.426926426427u,0 4555.336086586587u,0 4555.337086586587u,1.5 4556.3136266266265u,1.5 4556.314626626627u,0 4562.178866866867u,0 4562.179866866867u,1.5 4563.156406906906u,1.5 4563.1574069069065u,0 4565.111486986987u,0 4565.112486986987u,1.5 4569.021647147147u,1.5 4569.022647147147u,0 4569.999187187187u,0 4570.000187187187u,1.5 4576.841967467468u,1.5 4576.842967467468u,0 4577.819507507507u,0 4577.8205075075075u,1.5 4578.797047547547u,1.5 4578.798047547547u,0 4583.684747747748u,0 4583.685747747748u,1.5 4585.6398278278275u,1.5 4585.640827827828u,0 4586.617367867868u,0 4586.618367867868u,1.5 4587.594907907907u,1.5 4587.5959079079075u,0 4588.572447947948u,0 4588.573447947948u,1.5 4590.5275280280275u,1.5 4590.528528028028u,0 4591.505068068068u,0 4591.506068068068u,1.5 4597.370308308308u,1.5 4597.3713083083085u,0 4600.3029284284285u,0 4600.303928428429u,1.5 4601.280468468469u,1.5 4601.281468468469u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4607.145708708708u,1.5 4607.1467087087085u,0 4608.123248748749u,0 4608.124248748749u,1.5 4613.988488988989u,1.5 4613.989488988989u,0 4614.9660290290285u,0 4614.967029029029u,1.5 4615.943569069069u,1.5 4615.944569069069u,0 4616.921109109109u,0 4616.922109109109u,1.5 4617.898649149149u,1.5 4617.899649149149u,0 4620.83126926927u,0 4620.83226926927u,1.5 4622.786349349349u,1.5 4622.787349349349u,0 4623.763889389389u,0 4623.764889389389u,1.5 4627.674049549549u,1.5 4627.675049549549u,0 4629.6291296296295u,0 4629.63012962963u,1.5 4630.60666966967u,1.5 4630.60766966967u,0 4633.53928978979u,0 4633.54028978979u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4637.44944994995u,0 4637.45044994995u,1.5 4640.38207007007u,1.5 4640.38307007007u,0 4641.35961011011u,0 4641.36061011011u,1.5 4643.31469019019u,1.5 4643.31569019019u,0 4645.269770270271u,0 4645.270770270271u,1.5 4646.24731031031u,1.5 4646.24831031031u,0 4649.17993043043u,0 4649.180930430431u,1.5 4651.13501051051u,1.5 4651.1360105105105u,0 4652.11255055055u,0 4652.11355055055u,1.5 4653.090090590591u,1.5 4653.091090590591u,0 4654.06763063063u,0 4654.068630630631u,1.5 4655.045170670671u,1.5 4655.046170670671u,0 4657.000250750751u,0 4657.001250750751u,1.5 4657.977790790791u,1.5 4657.978790790791u,0 4658.9553308308305u,0 4658.956330830831u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4665.798111111111u,1.5 4665.799111111111u,0 4669.708271271272u,0 4669.709271271272u,1.5 4670.685811311311u,1.5 4670.686811311311u,0 4671.663351351351u,0 4671.664351351351u,1.5 4680.461211711711u,1.5 4680.4622117117115u,0 4682.416291791792u,0 4682.417291791792u,1.5 4683.393831831831u,1.5 4683.394831831832u,0 4685.348911911911u,0 4685.3499119119115u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4687.303991991992u,0 4687.304991991992u,1.5 4688.2815320320315u,1.5 4688.282532032032u,0 4689.259072072072u,0 4689.260072072072u,1.5 4691.214152152152u,1.5 4691.215152152152u,0 4692.191692192192u,0 4692.192692192192u,1.5 4693.1692322322315u,1.5 4693.170232232232u,0 4697.079392392392u,0 4697.080392392392u,1.5 4698.056932432432u,1.5 4698.057932432433u,0 4699.034472472473u,0 4699.035472472473u,1.5 4700.012012512512u,1.5 4700.013012512512u,0 4700.989552552552u,0 4700.990552552552u,1.5 4702.944632632632u,1.5 4702.945632632633u,0 4704.899712712712u,0 4704.900712712712u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4709.787412912912u,0 4709.7884129129125u,1.5 4713.697573073073u,1.5 4713.698573073073u,0 4718.585273273274u,0 4718.586273273274u,1.5 4720.540353353353u,1.5 4720.541353353353u,0 4722.495433433433u,0 4722.496433433434u,1.5 4725.428053553553u,1.5 4725.429053553553u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4734.225913913913u,1.5 4734.226913913913u,0 4735.203453953954u,0 4735.204453953954u,1.5 4736.180993993994u,1.5 4736.181993993994u,0 4740.091154154154u,0 4740.092154154154u,1.5 4744.001314314314u,1.5 4744.002314314314u,0 4744.978854354354u,0 4744.979854354354u,1.5 4745.956394394394u,1.5 4745.957394394394u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 4753.776714714714u,1.5 4753.777714714714u,0 4754.7542547547555u,0 4754.755254754756u,1.5 4755.731794794795u,1.5 4755.732794794795u,0 4756.709334834834u,0 4756.710334834835u,1.5 4757.686874874875u,1.5 4757.687874874875u,0 4760.619494994995u,0 4760.620494994995u,1.5 4761.597035035034u,1.5 4761.598035035035u,0 4763.552115115115u,0 4763.553115115115u,1.5 4767.462275275276u,1.5 4767.463275275276u,0 4770.394895395395u,0 4770.395895395395u,1.5 4772.349975475476u,1.5 4772.350975475476u,0 4774.305055555556u,0 4774.306055555556u,1.5 4778.215215715715u,1.5 4778.216215715715u,0 4781.147835835835u,0 4781.148835835836u,1.5 4784.0804559559565u,1.5 4784.081455955957u,0 4786.035536036035u,0 4786.036536036036u,1.5 4787.990616116116u,1.5 4787.991616116116u,0 4792.878316316316u,0 4792.879316316316u,1.5 4794.833396396396u,1.5 4794.834396396396u,0 4797.766016516516u,0 4797.767016516516u,1.5 4799.721096596597u,1.5 4799.722096596597u,0 4804.608796796797u,0 4804.609796796797u,1.5 4809.496496996997u,1.5 4809.497496996997u,0 4810.474037037036u,0 4810.475037037037u,1.5 4811.451577077077u,1.5 4811.452577077077u,0 4815.361737237236u,0 4815.362737237237u,1.5 4816.339277277278u,1.5 4816.340277277278u,0 4817.316817317317u,0 4817.317817317317u,1.5 4819.271897397397u,1.5 4819.272897397397u,0 4822.204517517517u,0 4822.205517517517u,1.5 4824.159597597598u,1.5 4824.160597597598u,0 4825.137137637637u,0 4825.138137637638u,1.5 4826.114677677678u,1.5 4826.115677677678u,0 4827.092217717717u,0 4827.093217717717u,1.5 4831.002377877878u,1.5 4831.003377877878u,0 4831.979917917918u,0 4831.980917917918u,1.5 4832.9574579579585u,1.5 4832.958457957959u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4843.710398398398u,1.5 4843.711398398398u,0 4844.687938438438u,0 4844.6889384384385u,1.5 4845.665478478479u,1.5 4845.666478478479u,0 4849.575638638638u,0 4849.5766386386385u,1.5 4850.553178678679u,1.5 4850.554178678679u,0 4851.530718718718u,0 4851.531718718718u,1.5 4852.508258758759u,1.5 4852.50925875876u,0 4853.485798798799u,0 4853.486798798799u,1.5 4854.463338838838u,1.5 4854.464338838839u,0 4855.440878878879u,0 4855.441878878879u,1.5 4857.395958958959u,1.5 4857.39695895896u,0 4865.21627927928u,0 4865.21727927928u,1.5 4870.10397947948u,1.5 4870.10497947948u,0 4872.0590595595595u,0 4872.06005955956u,1.5 4873.0365995996u,1.5 4873.0375995996u,0 4876.94675975976u,0 4876.947759759761u,1.5 4877.9242997998u,1.5 4877.9252997998u,0 4878.901839839839u,0 4878.9028398398395u,1.5 4879.87937987988u,1.5 4879.88037987988u,0 4880.85691991992u,0 4880.85791991992u,1.5 4881.83445995996u,1.5 4881.835459959961u,0 4885.74462012012u,0 4885.74562012012u,1.5 4886.7221601601605u,1.5 4886.723160160161u,0 4890.63232032032u,0 4890.63332032032u,1.5 4891.6098603603605u,1.5 4891.610860360361u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4895.52002052052u,1.5 4895.52102052052u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4903.34034084084u,1.5 4903.3413408408405u,0 4905.295420920921u,0 4905.296420920921u,1.5 4906.272960960961u,1.5 4906.273960960962u,0 4907.250501001001u,0 4907.251501001001u,1.5 4908.22804104104u,1.5 4908.229041041041u,0 4911.160661161161u,0 4911.161661161162u,1.5 4912.138201201201u,1.5 4912.139201201201u,0 4914.093281281282u,0 4914.094281281282u,1.5 4917.025901401401u,1.5 4917.026901401401u,0 4918.980981481482u,0 4918.981981481482u,1.5 4919.958521521521u,1.5 4919.959521521521u,0 4920.9360615615615u,0 4920.937061561562u,1.5 4921.913601601602u,1.5 4921.914601601602u,0 4923.868681681682u,0 4923.869681681682u,1.5 4924.846221721721u,1.5 4924.847221721721u,0 4930.711461961962u,0 4930.712461961963u,1.5 4931.689002002002u,1.5 4931.690002002002u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4935.599162162162u,0 4935.600162162163u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4939.509322322322u,1.5 4939.510322322322u,0 4940.486862362362u,0 4940.487862362363u,1.5 4945.3745625625625u,1.5 4945.375562562563u,0 4946.352102602603u,0 4946.353102602603u,1.5 4950.262262762763u,1.5 4950.263262762764u,0 4956.127503003003u,0 4956.128503003003u,1.5 4957.105043043042u,1.5 4957.1060430430425u,0 4964.925363363363u,0 4964.926363363364u,1.5 4965.902903403403u,1.5 4965.903903403403u,0 4969.813063563563u,0 4969.814063563564u,1.5 4970.790603603604u,1.5 4970.791603603604u,0 4971.768143643643u,0 4971.7691436436435u,1.5 4972.745683683684u,1.5 4972.746683683684u,0 4973.723223723723u,0 4973.724223723723u,1.5 4974.700763763764u,1.5 4974.701763763765u,0 4976.655843843843u,0 4976.6568438438435u,1.5 4977.633383883884u,1.5 4977.634383883884u,0 4978.610923923924u,0 4978.611923923924u,1.5 4983.498624124124u,1.5 4983.499624124124u,0 4984.476164164164u,0 4984.477164164165u,1.5 4985.453704204204u,1.5 4985.454704204204u,0 4986.431244244243u,0 4986.4322442442435u,1.5 4988.386324324324u,1.5 4988.387324324324u,0 4989.363864364364u,0 4989.364864364365u,1.5 4999.139264764765u,1.5 4999.140264764766u,0 5000.116804804805u,0 5000.117804804805u,1.5 5003.049424924925u,1.5 5003.050424924925u,0 5005.004505005005u,0 5005.005505005005u,1.5 5005.982045045044u,1.5 5005.9830450450445u,0 5007.937125125125u,0 5007.938125125125u,1.5 5014.779905405405u,1.5 5014.780905405405u,0 5016.734985485486u,0 5016.735985485486u,1.5 5017.712525525525u,1.5 5017.713525525525u,0 5018.690065565565u,0 5018.691065565566u,1.5 5020.645145645645u,1.5 5020.646145645645u,0 5024.555305805806u,0 5024.556305805806u,1.5 5025.532845845845u,1.5 5025.5338458458455u,0 5026.510385885886u,0 5026.511385885886u,1.5 5028.465465965966u,1.5 5028.466465965967u,0 5029.443006006006u,0 5029.444006006006u,1.5 5031.398086086087u,1.5 5031.399086086087u,0 5033.353166166166u,0 5033.354166166167u,1.5 5034.330706206206u,1.5 5034.331706206206u,0 5042.151026526526u,0 5042.152026526526u,1.5 5043.128566566566u,1.5 5043.129566566567u,0 5044.106106606607u,0 5044.107106606607u,1.5 5045.083646646646u,1.5 5045.084646646646u,0 5048.993806806807u,0 5048.994806806807u,1.5 5049.971346846846u,1.5 5049.972346846846u,0 5050.948886886887u,0 5050.949886886887u,1.5 5052.903966966967u,1.5 5052.904966966968u,0 5053.881507007007u,0 5053.882507007007u,1.5 5054.859047047046u,1.5 5054.8600470470465u,0 5057.791667167167u,0 5057.792667167168u,1.5 5059.746747247247u,1.5 5059.747747247247u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5067.567067567567u,0 5067.568067567568u,1.5 5068.544607607608u,1.5 5068.545607607608u,0 5071.477227727727u,0 5071.478227727727u,1.5 5072.454767767768u,1.5 5072.4557677677685u,0 5074.409847847847u,0 5074.410847847847u,1.5 5075.387387887888u,1.5 5075.388387887888u,0 5077.342467967968u,0 5077.3434679679685u,1.5 5078.320008008008u,1.5 5078.321008008008u,0 5079.297548048047u,0 5079.298548048047u,1.5 5081.252628128128u,1.5 5081.253628128128u,0 5082.230168168168u,0 5082.231168168169u,1.5 5084.185248248248u,1.5 5084.186248248248u,0 5085.1627882882885u,0 5085.163788288289u,1.5 5087.117868368368u,1.5 5087.118868368369u,0 5088.095408408408u,0 5088.096408408408u,1.5 5089.072948448448u,1.5 5089.073948448448u,0 5092.983108608609u,0 5092.984108608609u,1.5 5103.736049049048u,1.5 5103.737049049048u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5108.623749249249u,1.5 5108.624749249249u,0 5113.511449449449u,0 5113.512449449449u,1.5 5116.444069569569u,1.5 5116.44506956957u,0 5118.399149649649u,0 5118.400149649649u,1.5 5121.33176976977u,1.5 5121.3327697697705u,0 5122.30930980981u,0 5122.31030980981u,1.5 5123.286849849849u,1.5 5123.287849849849u,0 5129.1520900900905u,0 5129.153090090091u,1.5 5131.10717017017u,1.5 5131.1081701701705u,0 5132.08471021021u,0 5132.08571021021u,1.5 5134.0397902902905u,1.5 5134.040790290291u,0 5135.01733033033u,0 5135.01833033033u,1.5 5138.9274904904905u,1.5 5138.928490490491u,0 5141.860110610611u,0 5141.861110610611u,1.5 5142.83765065065u,1.5 5142.83865065065u,0 5143.8151906906905u,0 5143.816190690691u,1.5 5148.702890890891u,1.5 5148.703890890891u,0 5154.568131131131u,0 5154.569131131131u,1.5 5155.545671171171u,1.5 5155.5466711711715u,0 5156.523211211211u,0 5156.524211211211u,1.5 5157.500751251251u,1.5 5157.501751251251u,0 5159.455831331331u,0 5159.456831331331u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5163.3659914914915u,0 5163.366991491492u,1.5 5164.343531531531u,1.5 5164.344531531531u,0 5167.276151651651u,0 5167.277151651651u,1.5 5169.231231731731u,1.5 5169.232231731731u,0 5170.208771771772u,0 5170.2097717717725u,1.5 5173.1413918918915u,1.5 5173.142391891892u,0 5174.118931931932u,0 5174.119931931932u,1.5 5175.096471971972u,1.5 5175.0974719719725u,0 5180.961712212212u,0 5180.962712212212u,1.5 5181.939252252252u,1.5 5181.940252252252u,0 5182.9167922922925u,0 5182.917792292293u,1.5 5185.849412412412u,1.5 5185.850412412412u,0 5186.826952452452u,0 5186.827952452452u,1.5 5187.8044924924925u,1.5 5187.805492492493u,0 5189.759572572572u,0 5189.7605725725725u,1.5 5190.737112612613u,1.5 5190.738112612613u,0 5191.714652652652u,0 5191.715652652652u,1.5 5193.669732732732u,1.5 5193.670732732732u,0 5194.647272772773u,0 5194.648272772773u,1.5 5197.5798928928925u,1.5 5197.580892892893u,0 5203.445133133133u,0 5203.446133133133u,1.5 5207.3552932932935u,1.5 5207.356293293294u,0 5208.332833333333u,0 5208.333833333333u,1.5 5211.265453453453u,1.5 5211.266453453453u,0 5213.220533533533u,0 5213.221533533533u,1.5 5214.198073573573u,1.5 5214.1990735735735u,0 5216.153153653653u,0 5216.154153653653u,1.5 5217.1306936936935u,1.5 5217.131693693694u,0 5218.108233733733u,0 5218.109233733733u,1.5 5219.085773773774u,1.5 5219.086773773774u,0 5220.063313813814u,0 5220.064313813814u,1.5 5221.040853853853u,1.5 5221.041853853853u,0 5223.973473973974u,0 5223.974473973974u,1.5 5224.951014014014u,1.5 5224.952014014014u,0 5225.928554054053u,0 5225.929554054053u,1.5 5228.861174174174u,1.5 5228.8621741741745u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5235.703954454454u,0 5235.704954454454u,1.5 5239.614114614615u,1.5 5239.615114614615u,0 5244.501814814815u,0 5244.502814814815u,1.5 5245.479354854854u,1.5 5245.480354854854u,0 5246.4568948948945u,0 5246.457894894895u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5258.187375375375u,0 5258.1883753753755u,1.5 5259.164915415415u,1.5 5259.165915415415u,0 5261.1199954954955u,0 5261.120995495496u,1.5 5262.097535535535u,1.5 5262.098535535535u,0 5263.075075575575u,0 5263.0760755755755u,1.5 5266.0076956956955u,1.5 5266.008695695696u,0 5266.985235735735u,0 5266.986235735735u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5274.805556056056u,0 5274.806556056056u,1.5 5281.648336336336u,1.5 5281.649336336336u,0 5282.625876376376u,0 5282.6268763763765u,1.5 5284.580956456457u,1.5 5284.581956456457u,0 5288.491116616617u,0 5288.492116616617u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5297.288976976977u,0 5297.289976976977u,1.5 5300.221597097097u,1.5 5300.222597097098u,0 5301.199137137137u,0 5301.200137137137u,1.5 5303.154217217217u,1.5 5303.155217217217u,0 5309.019457457458u,0 5309.020457457458u,1.5 5310.974537537537u,1.5 5310.975537537537u,0 5311.952077577577u,0 5311.9530775775775u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5316.839777777778u,1.5 5316.840777777778u,0 5319.7723978978975u,0 5319.773397897898u,1.5 5327.592718218218u,1.5 5327.593718218218u,0 5331.502878378378u,0 5331.503878378378u,1.5 5332.480418418419u,1.5 5332.481418418419u,0 5333.457958458459u,0 5333.458958458459u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5344.210898898898u,0 5344.211898898899u,1.5 5345.188438938939u,1.5 5345.189438938939u,0 5347.143519019019u,0 5347.144519019019u,1.5 5348.121059059059u,1.5 5348.122059059059u,0 5350.076139139139u,0 5350.077139139139u,1.5 5352.031219219219u,1.5 5352.032219219219u,0 5357.89645945946u,0 5357.89745945946u,1.5 5359.851539539539u,1.5 5359.852539539539u,0 5360.829079579579u,0 5360.830079579579u,1.5 5365.71677977978u,1.5 5365.71777977978u,0 5369.62693993994u,0 5369.62793993994u,1.5 5370.60447997998u,1.5 5370.60547997998u,0 5371.58202002002u,0 5371.58302002002u,1.5 5376.46972022022u,1.5 5376.47072022022u,0 5377.447260260261u,0 5377.448260260261u,1.5 5378.4248003003u,1.5 5378.425800300301u,0 5380.37988038038u,0 5380.38088038038u,1.5 5382.334960460461u,1.5 5382.335960460461u,0 5387.222660660661u,0 5387.223660660661u,1.5 5392.110360860861u,1.5 5392.111360860861u,0 5393.0879009009u,0 5393.088900900901u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5400.908221221221u,0 5400.909221221221u,1.5 5401.885761261262u,1.5 5401.886761261262u,0 5404.818381381381u,0 5404.819381381381u,1.5 5408.728541541541u,1.5 5408.729541541541u,0 5409.706081581581u,0 5409.707081581581u,1.5 5411.661161661662u,1.5 5411.662161661662u,0 5412.638701701701u,0 5412.639701701702u,1.5 5415.571321821822u,1.5 5415.572321821822u,0 5417.526401901901u,0 5417.527401901902u,1.5 5418.503941941942u,1.5 5418.504941941942u,0 5421.436562062062u,0 5421.437562062062u,1.5 5422.414102102102u,1.5 5422.4151021021025u,0 5423.391642142142u,0 5423.392642142142u,1.5 5424.369182182182u,1.5 5424.370182182182u,0 5425.346722222222u,0 5425.347722222222u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5434.144582582582u,0 5434.145582582582u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5442.942442942943u,0 5442.943442942943u,1.5 5444.897523023023u,1.5 5444.898523023023u,0 5446.852603103103u,0 5446.8536031031035u,1.5 5447.830143143143u,1.5 5447.831143143143u,0 5448.807683183183u,0 5448.808683183183u,1.5 5450.762763263264u,1.5 5450.763763263264u,0 5452.717843343343u,0 5452.718843343343u,1.5 5456.628003503503u,1.5 5456.629003503504u,0 5458.583083583583u,0 5458.584083583583u,1.5 5459.5606236236235u,1.5 5459.561623623624u,0 5461.515703703703u,0 5461.516703703704u,1.5 5466.403403903903u,1.5 5466.404403903904u,0 5467.380943943944u,0 5467.381943943944u,1.5 5468.358483983984u,1.5 5468.359483983984u,0 5469.336024024024u,0 5469.337024024024u,1.5 5471.291104104104u,1.5 5471.2921041041045u,0 5473.246184184184u,0 5473.247184184184u,1.5 5474.223724224224u,1.5 5474.224724224224u,0 5475.201264264265u,0 5475.202264264265u,1.5 5476.178804304304u,1.5 5476.1798043043045u,0 5478.133884384384u,0 5478.134884384384u,1.5 5479.1114244244245u,1.5 5479.112424424425u,0 5481.066504504504u,0 5481.0675045045045u,1.5 5482.044044544544u,1.5 5482.045044544544u,0 5483.9991246246245u,0 5484.000124624625u,1.5 5484.976664664665u,1.5 5484.977664664665u,0 5490.841904904904u,0 5490.842904904905u,1.5 5491.819444944945u,1.5 5491.820444944945u,0 5492.796984984985u,0 5492.797984984985u,1.5 5495.729605105105u,1.5 5495.7306051051055u,0 5497.684685185185u,0 5497.685685185185u,1.5 5498.662225225225u,1.5 5498.663225225225u,0 5503.5499254254255u,0 5503.550925425426u,1.5 5504.527465465466u,1.5 5504.528465465466u,0 5511.370245745745u,0 5511.371245745745u,1.5 5513.3253258258255u,1.5 5513.326325825826u,0 5520.168106106106u,0 5520.1691061061065u,1.5 5522.123186186186u,1.5 5522.124186186186u,0 5524.078266266267u,0 5524.079266266267u,1.5 5525.055806306306u,1.5 5525.0568063063065u,0 5527.9884264264265u,0 5527.989426426427u,1.5 5528.965966466467u,1.5 5528.966966466467u,0 5529.943506506506u,0 5529.9445065065065u,1.5 5533.853666666667u,1.5 5533.854666666667u,0 5534.831206706706u,0 5534.8322067067065u,1.5 5539.718906906906u,1.5 5539.7199069069065u,0 5544.606607107107u,0 5544.6076071071075u,1.5 5547.539227227227u,1.5 5547.540227227227u,0 5548.516767267268u,0 5548.517767267268u,1.5 5551.449387387387u,1.5 5551.450387387387u,0 5553.404467467468u,0 5553.405467467468u,1.5 5554.382007507507u,1.5 5554.3830075075075u,0 5557.3146276276275u,0 5557.315627627628u,1.5 5559.269707707707u,1.5 5559.2707077077075u,0 5564.157407907907u,0 5564.1584079079075u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5569.045108108108u,0 5569.0461081081085u,1.5 5574.910348348348u,1.5 5574.911348348348u,0 5575.887888388388u,0 5575.888888388388u,1.5 5578.820508508508u,1.5 5578.8215085085085u,0 5584.685748748749u,0 5584.686748748749u,1.5 5585.663288788789u,1.5 5585.664288788789u,0 5587.618368868869u,0 5587.619368868869u,1.5 5596.4162292292285u,1.5 5596.417229229229u,0 5598.371309309309u,0 5598.3723093093095u,1.5 5600.326389389389u,1.5 5600.327389389389u,0 5601.303929429429u,0 5601.30492942943u,1.5 5602.28146946947u,1.5 5602.28246946947u,0 5604.236549549549u,0 5604.237549549549u,1.5 5606.1916296296295u,1.5 5606.19262962963u,0 5607.16916966967u,0 5607.17016966967u,1.5 5608.146709709709u,1.5 5608.1477097097095u,0 5609.12424974975u,0 5609.12524974975u,1.5 5614.01194994995u,1.5 5614.01294994995u,0 5614.98948998999u,0 5614.99048998999u,1.5 5615.9670300300295u,1.5 5615.96803003003u,0 5616.94457007007u,0 5616.94557007007u,1.5 5618.89965015015u,1.5 5618.90065015015u,0 5619.87719019019u,0 5619.87819019019u,1.5 5620.8547302302295u,1.5 5620.85573023023u,0 5623.78735035035u,0 5623.78835035035u,1.5 5626.719970470471u,1.5 5626.720970470471u,0 5627.69751051051u,0 5627.6985105105105u,1.5 5628.67505055055u,1.5 5628.67605055055u,0 5630.63013063063u,0 5630.631130630631u,1.5 5631.607670670671u,1.5 5631.608670670671u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5641.383071071071u,1.5 5641.384071071071u,0 5642.360611111111u,0 5642.361611111111u,1.5 5643.338151151151u,1.5 5643.339151151151u,0 5644.315691191191u,0 5644.316691191191u,1.5 5645.2932312312305u,1.5 5645.294231231231u,0 5647.248311311311u,0 5647.249311311311u,1.5 5650.180931431431u,1.5 5650.181931431432u,0 5652.136011511511u,0 5652.137011511511u,1.5 5656.046171671672u,1.5 5656.047171671672u,0 5657.023711711711u,0 5657.0247117117115u,1.5 5658.001251751752u,1.5 5658.002251751752u,0 5659.956331831831u,0 5659.957331831832u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5662.888951951952u,0 5662.889951951952u,1.5 5668.754192192192u,1.5 5668.755192192192u,0 5672.664352352352u,0 5672.665352352352u,1.5 5674.619432432432u,1.5 5674.620432432433u,0 5675.596972472473u,0 5675.597972472473u,1.5 5680.484672672673u,1.5 5680.485672672673u,0 5685.372372872873u,0 5685.373372872873u,1.5 5686.349912912912u,1.5 5686.3509129129125u,0 5687.327452952953u,0 5687.328452952953u,1.5 5692.215153153153u,1.5 5692.216153153153u,0 5693.192693193193u,0 5693.193693193193u,1.5 5694.1702332332325u,1.5 5694.171233233233u,0 5696.125313313313u,0 5696.126313313313u,1.5 5698.080393393393u,1.5 5698.081393393393u,0 5700.035473473474u,0 5700.036473473474u,1.5 5701.990553553553u,1.5 5701.991553553553u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5712.743493993994u,1.5 5712.744493993994u,0 5713.721034034033u,0 5713.722034034034u,1.5 5714.698574074074u,1.5 5714.699574074074u,0 5719.586274274275u,0 5719.587274274275u,1.5 5721.541354354354u,1.5 5721.542354354354u,0 5722.518894394394u,0 5722.519894394394u,1.5 5723.496434434434u,1.5 5723.497434434435u,0 5724.473974474475u,0 5724.474974474475u,1.5 5725.451514514514u,1.5 5725.452514514514u,0 5728.384134634634u,0 5728.385134634635u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5731.316754754755u,1.5 5731.317754754755u,0 5732.294294794795u,0 5732.295294794795u,1.5 5735.226914914914u,1.5 5735.227914914914u,0 5736.204454954955u,0 5736.205454954955u,1.5 5737.181994994995u,1.5 5737.182994994995u,0 5739.137075075075u,0 5739.138075075075u,1.5 5740.114615115115u,1.5 5740.115615115115u,0 5741.092155155155u,0 5741.093155155155u,1.5 5745.002315315315u,1.5 5745.003315315315u,0 5750.867555555555u,0 5750.868555555555u,1.5 5753.800175675676u,1.5 5753.801175675676u,0 5760.6429559559565u,0 5760.643955955957u,1.5 5762.598036036035u,1.5 5762.599036036036u,0 5763.575576076076u,0 5763.576576076076u,1.5 5766.508196196196u,1.5 5766.509196196196u,0 5767.485736236235u,0 5767.486736236236u,1.5 5768.463276276277u,1.5 5768.464276276277u,0 5769.440816316316u,0 5769.441816316316u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5775.3060565565565u,1.5 5775.307056556557u,0 5776.283596596597u,0 5776.284596596597u,1.5 5777.261136636636u,1.5 5777.262136636637u,0 5778.238676676677u,0 5778.239676676677u,1.5 5779.216216716716u,1.5 5779.217216716716u,0 5780.1937567567575u,0 5780.194756756758u,1.5 5781.171296796797u,1.5 5781.172296796797u,0 5782.148836836836u,0 5782.149836836837u,1.5 5785.0814569569575u,1.5 5785.082456956958u,0 5791.924237237236u,0 5791.925237237237u,1.5 5794.8568573573575u,1.5 5794.857857357358u,0 5795.834397397397u,0 5795.835397397397u,1.5 5796.811937437437u,1.5 5796.8129374374375u,0 5797.789477477478u,0 5797.790477477478u,1.5 5798.767017517517u,1.5 5798.768017517517u,0 5802.677177677678u,0 5802.678177677678u,1.5 5803.654717717717u,1.5 5803.655717717717u,0 5804.632257757758u,0 5804.633257757759u,1.5 5806.587337837837u,1.5 5806.588337837838u,0 5807.564877877878u,0 5807.565877877878u,1.5 5809.5199579579585u,1.5 5809.520957957959u,0 5811.475038038037u,0 5811.476038038038u,1.5 5812.452578078078u,1.5 5812.453578078078u,0 5814.4076581581585u,0 5814.408658158159u,1.5 5816.362738238237u,1.5 5816.363738238238u,0 5818.317818318318u,0 5818.318818318318u,1.5 5820.272898398398u,1.5 5820.273898398398u,0 5821.250438438438u,0 5821.2514384384385u,1.5 5822.227978478479u,1.5 5822.228978478479u,0 5827.115678678679u,0 5827.116678678679u,1.5 5834.935998998999u,1.5 5834.936998998999u,0 5836.891079079079u,0 5836.892079079079u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5839.823699199199u,0 5839.824699199199u,1.5 5842.756319319319u,1.5 5842.757319319319u,0 5843.7338593593595u,0 5843.73485935936u,1.5 5845.688939439439u,1.5 5845.6899394394395u,0 5846.66647947948u,0 5846.66747947948u,1.5 5847.644019519519u,1.5 5847.645019519519u,0 5849.5990995996u,0 5849.6000995996u,1.5 5850.576639639639u,1.5 5850.5776396396395u,0 5851.55417967968u,0 5851.55517967968u,1.5 5857.41941991992u,1.5 5857.42041991992u,0 5858.39695995996u,0 5858.397959959961u,1.5 5859.3745u,1.5 5859.3755u,0 5860.352040040039u,0 5860.35304004004u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5863.2846601601605u,0 5863.285660160161u,1.5 5864.2622002002u,1.5 5864.2632002002u,0 5865.239740240239u,0 5865.24074024024u,1.5 5866.217280280281u,1.5 5866.218280280281u,0 5867.19482032032u,0 5867.19582032032u,1.5 5871.104980480481u,1.5 5871.105980480481u,0 5872.08252052052u,0 5872.08352052052u,1.5 5873.0600605605605u,1.5 5873.061060560561u,0 5877.947760760761u,0 5877.948760760762u,1.5 5878.925300800801u,1.5 5878.926300800801u,0 5879.90284084084u,0 5879.9038408408405u,1.5 5880.880380880881u,1.5 5880.881380880881u,0 5881.857920920921u,0 5881.858920920921u,1.5 5882.835460960961u,1.5 5882.836460960962u,0 5883.813001001001u,0 5883.814001001001u,1.5 5885.768081081081u,1.5 5885.769081081081u,0 5888.700701201201u,0 5888.701701201201u,1.5 5889.67824124124u,1.5 5889.679241241241u,0 5891.633321321321u,0 5891.634321321321u,1.5 5892.6108613613615u,1.5 5892.611861361362u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5896.521021521521u,1.5 5896.522021521521u,0 5897.4985615615615u,0 5897.499561561562u,1.5 5899.453641641641u,1.5 5899.4546416416415u,0 5900.431181681682u,0 5900.432181681682u,1.5 5901.408721721721u,1.5 5901.409721721721u,0 5902.386261761762u,0 5902.387261761763u,1.5 5903.363801801802u,1.5 5903.364801801802u,0 5904.341341841841u,0 5904.3423418418415u,1.5 5905.318881881882u,1.5 5905.319881881882u,0 5907.273961961962u,0 5907.274961961963u,1.5 5908.251502002002u,1.5 5908.252502002002u,0 5910.206582082082u,0 5910.207582082082u,1.5 5911.184122122122u,1.5 5911.185122122122u,0 5913.139202202202u,0 5913.140202202202u,1.5 5921.9370625625625u,1.5 5921.938062562563u,0 5922.914602602603u,0 5922.915602602603u,1.5 5923.892142642642u,1.5 5923.8931426426425u,0 5926.824762762763u,0 5926.825762762764u,1.5 5927.802302802803u,1.5 5927.803302802803u,0 5930.734922922923u,0 5930.735922922923u,1.5 5931.712462962963u,1.5 5931.713462962964u,0 5935.622623123123u,0 5935.623623123123u,1.5 5942.465403403403u,1.5 5942.466403403403u,0 5944.420483483484u,0 5944.421483483484u,1.5 5945.398023523523u,1.5 5945.399023523523u,0 5946.375563563563u,0 5946.376563563564u,1.5 5949.308183683684u,1.5 5949.309183683684u,0 5950.285723723723u,0 5950.286723723723u,1.5 5952.240803803804u,1.5 5952.241803803804u,0 5953.218343843843u,0 5953.2193438438435u,1.5 5954.195883883884u,1.5 5954.196883883884u,0 5958.106044044043u,0 5958.1070440440435u,1.5 5959.083584084084u,1.5 5959.084584084084u,0 5962.993744244243u,0 5962.9947442442435u,1.5 5963.971284284285u,1.5 5963.972284284285u,0 5964.948824324324u,0 5964.949824324324u,1.5 5965.926364364364u,1.5 5965.927364364365u,0 5967.881444444444u,0 5967.882444444444u,1.5 5968.858984484485u,1.5 5968.859984484485u,0 5970.814064564564u,0 5970.815064564565u,1.5 5971.791604604605u,1.5 5971.792604604605u,0 5972.769144644644u,0 5972.7701446446445u,1.5 5973.746684684685u,1.5 5973.747684684685u,0 5974.724224724724u,0 5974.725224724724u,1.5 5976.679304804805u,1.5 5976.680304804805u,0 5977.656844844844u,0 5977.6578448448445u,1.5 5980.589464964965u,1.5 5980.590464964966u,0 5981.567005005005u,0 5981.568005005005u,1.5 5992.319945445445u,1.5 5992.320945445445u,0 5993.297485485486u,0 5993.298485485486u,1.5 5994.275025525525u,1.5 5994.276025525525u,0 5995.252565565565u,0 5995.253565565566u,1.5 5996.230105605606u,1.5 5996.231105605606u,0 5997.207645645645u,0 5997.208645645645u,1.5 6001.117805805806u,1.5 6001.118805805806u,0 6002.095345845845u,0 6002.0963458458455u,1.5 6013.825826326326u,1.5 6013.826826326326u,0 6014.803366366366u,0 6014.804366366367u,1.5 6019.691066566566u,1.5 6019.692066566567u,0 6020.668606606607u,0 6020.669606606607u,1.5 6024.578766766767u,1.5 6024.5797667667675u,0 6025.556306806807u,0 6025.557306806807u,1.5 6029.466466966967u,1.5 6029.467466966968u,0 6031.421547047046u,0 6031.4225470470465u,1.5 6035.331707207207u,1.5 6035.332707207207u,0 6036.309247247247u,0 6036.310247247247u,1.5 6038.264327327327u,1.5 6038.265327327327u,0 6045.107107607608u,0 6045.108107607608u,1.5 6046.084647647647u,1.5 6046.085647647647u,0 6048.039727727727u,0 6048.040727727727u,1.5 6049.017267767768u,1.5 6049.0182677677685u,0 6049.994807807808u,0 6049.995807807808u,1.5 6050.972347847847u,1.5 6050.973347847847u,0 6051.949887887888u,0 6051.950887887888u,1.5 6052.927427927928u,1.5 6052.928427927928u,0 6053.904967967968u,0 6053.9059679679685u,1.5 6061.7252882882885u,1.5 6061.726288288289u,0 6063.680368368368u,0 6063.681368368369u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6073.455768768769u,0 6073.4567687687695u,1.5 6077.365928928929u,1.5 6077.366928928929u,0 6078.343468968969u,0 6078.3444689689695u,1.5 6079.321009009009u,1.5 6079.322009009009u,0 6080.298549049048u,0 6080.299549049048u,1.5 6082.253629129129u,1.5 6082.254629129129u,0 6083.231169169169u,0 6083.2321691691695u,1.5 6084.208709209209u,1.5 6084.209709209209u,0 6085.186249249249u,0 6085.187249249249u,1.5 6087.141329329329u,1.5 6087.142329329329u,0 6088.118869369369u,0 6088.11986936937u,1.5 6090.073949449449u,1.5 6090.074949449449u,0 6091.0514894894895u,0 6091.05248948949u,1.5 6092.029029529529u,1.5 6092.030029529529u,0 6094.961649649649u,0 6094.962649649649u,1.5 6095.93918968969u,1.5 6095.94018968969u,0 6096.916729729729u,0 6096.917729729729u,1.5 6098.87180980981u,1.5 6098.87280980981u,0 6099.849349849849u,0 6099.850349849849u,1.5 6103.75951001001u,1.5 6103.76051001001u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6110.6022902902905u,0 6110.603290290291u,1.5 6111.57983033033u,1.5 6111.58083033033u,0 6114.51245045045u,0 6114.51345045045u,1.5 6116.46753053053u,1.5 6116.46853053053u,0 6117.44507057057u,0 6117.446070570571u,1.5 6120.3776906906905u,1.5 6120.378690690691u,0 6121.35523073073u,0 6121.35623073073u,1.5 6122.332770770771u,1.5 6122.3337707707715u,0 6123.310310810811u,0 6123.311310810811u,1.5 6124.28785085085u,1.5 6124.28885085085u,0 6128.198011011011u,0 6128.199011011011u,1.5 6129.17555105105u,1.5 6129.17655105105u,0 6130.1530910910915u,0 6130.154091091092u,1.5 6132.108171171171u,1.5 6132.1091711711715u,0 6134.063251251251u,0 6134.064251251251u,1.5 6136.995871371371u,1.5 6136.9968713713715u,0 6142.861111611612u,0 6142.862111611612u,1.5 6143.838651651651u,1.5 6143.839651651651u,0 6144.8161916916915u,0 6144.817191691692u,1.5 6147.748811811812u,1.5 6147.749811811812u,0 6148.726351851851u,0 6148.727351851851u,1.5 6149.7038918918915u,1.5 6149.704891891892u,0 6151.658971971972u,0 6151.6599719719725u,1.5 6152.636512012012u,1.5 6152.637512012012u,0 6156.546672172172u,0 6156.5476721721725u,1.5 6157.524212212212u,1.5 6157.525212212212u,0 6158.501752252252u,0 6158.502752252252u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6161.434372372372u,0 6161.4353723723725u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6163.389452452452u,0 6163.390452452452u,1.5 6164.3669924924925u,1.5 6164.367992492493u,0 6169.2546926926925u,0 6169.255692692693u,1.5 6170.232232732732u,1.5 6170.233232732732u,0 6171.209772772773u,0 6171.210772772773u,1.5 6172.187312812813u,1.5 6172.188312812813u,0 6173.164852852852u,0 6173.165852852852u,1.5 6175.119932932933u,1.5 6175.120932932933u,0 6180.985173173173u,0 6180.9861731731735u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6190.760573573573u,0 6190.7615735735735u,1.5 6195.648273773774u,1.5 6195.649273773774u,0 6196.625813813814u,0 6196.626813813814u,1.5 6197.603353853853u,1.5 6197.604353853853u,0 6202.491054054053u,0 6202.492054054053u,1.5 6207.378754254254u,1.5 6207.379754254254u,0 6213.2439944944945u,0 6213.244994494495u,1.5 6214.221534534534u,1.5 6214.222534534534u,0 6215.199074574574u,0 6215.2000745745745u,1.5 6217.154154654654u,1.5 6217.155154654654u,0 6219.109234734734u,0 6219.110234734734u,1.5 6220.086774774775u,1.5 6220.087774774775u,0 6223.0193948948945u,0 6223.020394894895u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6230.839715215215u,0 6230.840715215215u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6234.749875375375u,0 6234.7508753753755u,1.5 6238.660035535535u,1.5 6238.661035535535u,0 6239.637575575575u,0 6239.6385755755755u,1.5 6240.615115615616u,1.5 6240.616115615616u,0 6244.525275775776u,0 6244.526275775776u,1.5 6247.4578958958955u,1.5 6247.458895895896u,0 6250.390516016016u,0 6250.391516016016u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6253.323136136136u,0 6253.324136136136u,1.5 6255.278216216216u,1.5 6255.279216216216u,0 6256.255756256256u,0 6256.256756256256u,1.5 6257.233296296296u,1.5 6257.234296296297u,0 6258.210836336336u,0 6258.211836336336u,1.5 6259.188376376376u,1.5 6259.1893763763765u,0 6260.165916416417u,0 6260.166916416417u,1.5 6261.143456456457u,1.5 6261.144456456457u,0 6262.120996496496u,0 6262.121996496497u,1.5 6263.098536536536u,1.5 6263.099536536536u,0 6268.963776776777u,0 6268.964776776777u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6274.829017017017u,0 6274.830017017017u,1.5 6275.806557057057u,1.5 6275.807557057057u,0 6276.784097097097u,0 6276.785097097098u,1.5 6277.761637137137u,1.5 6277.762637137137u,0 6278.739177177177u,0 6278.740177177177u,1.5 6279.716717217217u,1.5 6279.717717217217u,0 6280.694257257258u,0 6280.695257257258u,1.5 6281.671797297297u,1.5 6281.672797297298u,0 6282.649337337337u,0 6282.650337337337u,1.5 6283.626877377377u,1.5 6283.627877377377u,0 6285.581957457458u,0 6285.582957457458u,1.5 6286.559497497497u,1.5 6286.560497497498u,0 6287.537037537537u,0 6287.538037537537u,1.5 6288.514577577577u,1.5 6288.5155775775775u,0 6290.469657657658u,0 6290.470657657658u,1.5 6293.402277777778u,1.5 6293.403277777778u,0 6296.3348978978975u,0 6296.335897897898u,1.5 6297.312437937938u,1.5 6297.313437937938u,0 6299.267518018018u,0 6299.268518018018u,1.5 6300.245058058058u,1.5 6300.246058058058u,0 6301.222598098098u,0 6301.223598098099u,1.5 6303.177678178178u,1.5 6303.178678178178u,0 6307.087838338338u,0 6307.088838338338u,1.5 6308.065378378378u,1.5 6308.066378378378u,0 6309.042918418419u,0 6309.043918418419u,1.5 6310.997998498498u,1.5 6310.998998498499u,0 6311.975538538538u,0 6311.976538538538u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6320.773398898898u,0 6320.774398898899u,1.5 6322.728478978979u,1.5 6322.729478978979u,0 6324.683559059059u,0 6324.684559059059u,1.5 6325.661099099099u,1.5 6325.6620990991u,0 6326.638639139139u,0 6326.639639139139u,1.5 6327.616179179179u,1.5 6327.617179179179u,0 6330.548799299299u,0 6330.5497992993u,1.5 6331.526339339339u,1.5 6331.527339339339u,0 6332.503879379379u,0 6332.504879379379u,1.5 6338.36911961962u,1.5 6338.37011961962u,0 6344.23435985986u,0 6344.23535985986u,1.5 6345.211899899899u,1.5 6345.2128998999u,0 6346.18943993994u,0 6346.19043993994u,1.5 6347.16697997998u,1.5 6347.16797997998u,0 6348.14452002002u,0 6348.14552002002u,1.5 6350.0996001001u,1.5 6350.100600100101u,0 6351.07714014014u,0 6351.07814014014u,1.5 6352.05468018018u,1.5 6352.05568018018u,0 6355.96484034034u,0 6355.96584034034u,1.5 6359.8750005005u,1.5 6359.876000500501u,0 6360.85254054054u,0 6360.85354054054u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6364.7627007007u,1.5 6364.763700700701u,0 6367.695320820821u,0 6367.696320820821u,1.5 6369.6504009009u,1.5 6369.651400900901u,0 6370.627940940941u,0 6370.628940940941u,1.5 6372.583021021021u,1.5 6372.584021021021u,0 6373.560561061061u,0 6373.561561061061u,1.5 6374.538101101101u,1.5 6374.539101101102u,0 6376.493181181181u,0 6376.494181181181u,1.5 6378.448261261262u,1.5 6378.449261261262u,0 6381.380881381381u,0 6381.381881381381u,1.5 6383.335961461462u,1.5 6383.336961461462u,0 6386.268581581581u,0 6386.269581581581u,1.5 6389.201201701701u,1.5 6389.202201701702u,0 6391.156281781782u,0 6391.157281781782u,1.5 6393.111361861862u,1.5 6393.112361861862u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6396.043981981982u,0 6396.044981981982u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6399.954142142142u,0 6399.955142142142u,1.5 6400.931682182182u,1.5 6400.932682182182u,0 6402.886762262263u,0 6402.887762262263u,1.5 6403.864302302302u,1.5 6403.865302302303u,0 6404.841842342342u,0 6404.842842342342u,1.5 6411.684622622623u,1.5 6411.685622622623u,0 6412.662162662663u,0 6412.663162662663u,1.5 6413.639702702702u,1.5 6413.640702702703u,0 6414.617242742742u,0 6414.618242742742u,1.5 6416.572322822823u,1.5 6416.573322822823u,0 6419.504942942943u,0 6419.505942942943u,1.5 6421.460023023023u,1.5 6421.461023023023u,0 6422.437563063063u,0 6422.438563063063u,1.5 6427.325263263264u,1.5 6427.326263263264u,0 6428.302803303303u,0 6428.3038033033035u,1.5 6432.212963463464u,1.5 6432.213963463464u,0 6433.190503503503u,0 6433.191503503504u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6436.1231236236235u,1.5 6436.124123623624u,0 6438.078203703703u,0 6438.079203703704u,1.5 6439.055743743743u,1.5 6439.056743743743u,0 6442.965903903903u,0 6442.966903903904u,1.5 6443.943443943944u,1.5 6443.944443943944u,0 6446.876064064064u,0 6446.877064064064u,1.5 6447.853604104104u,1.5 6447.8546041041045u,0 6448.831144144144u,0 6448.832144144144u,1.5 6449.808684184184u,1.5 6449.809684184184u,0 6450.786224224224u,0 6450.787224224224u,1.5 6451.763764264265u,1.5 6451.764764264265u,0 6452.741304304304u,0 6452.7423043043045u,1.5 6456.651464464465u,1.5 6456.652464464465u,0 6457.629004504504u,0 6457.6300045045045u,1.5 6460.5616246246245u,1.5 6460.562624624625u,0 6461.539164664665u,0 6461.540164664665u,1.5 6466.426864864865u,1.5 6466.427864864865u,0 6467.404404904904u,0 6467.405404904905u,1.5 6468.381944944945u,1.5 6468.382944944945u,0 6469.359484984985u,0 6469.360484984985u,1.5 6470.337025025025u,1.5 6470.338025025025u,0 6471.314565065065u,0 6471.315565065065u,1.5 6472.292105105105u,1.5 6472.2931051051055u,0 6473.269645145145u,0 6473.270645145145u,1.5 6474.247185185185u,1.5 6474.248185185185u,0 6477.179805305305u,0 6477.1808053053055u,1.5 6478.157345345345u,1.5 6478.158345345345u,0 6483.045045545545u,0 6483.046045545545u,1.5 6485.977665665666u,1.5 6485.978665665666u,0 6486.955205705705u,0 6486.9562057057055u,1.5 6487.932745745745u,1.5 6487.933745745745u,0 6489.8878258258255u,0 6489.888825825826u,1.5 6491.842905905905u,1.5 6491.843905905906u,0 6494.775526026026u,0 6494.776526026026u,1.5 6496.730606106106u,1.5 6496.7316061061065u,0 6500.640766266267u,0 6500.641766266267u,1.5 6501.618306306306u,1.5 6501.6193063063065u,0 6502.595846346346u,0 6502.596846346346u,1.5 6505.528466466467u,1.5 6505.529466466467u,0 6508.461086586587u,0 6508.462086586587u,1.5 6510.416166666667u,1.5 6510.417166666667u,0 6512.371246746747u,0 6512.372246746747u,1.5 6515.303866866867u,1.5 6515.304866866867u,0 6516.281406906906u,0 6516.2824069069065u,1.5 6517.258946946947u,1.5 6517.259946946947u,0 6519.2140270270265u,0 6519.215027027027u,1.5 6520.191567067067u,1.5 6520.192567067067u,0 6521.169107107107u,0 6521.1701071071075u,1.5 6522.146647147147u,1.5 6522.147647147147u,0 6523.124187187187u,0 6523.125187187187u,1.5 6524.101727227227u,1.5 6524.102727227227u,0 6525.079267267268u,0 6525.080267267268u,1.5 6526.056807307307u,1.5 6526.0578073073075u,0 6528.011887387387u,0 6528.012887387387u,1.5 6529.966967467468u,1.5 6529.967967467468u,0 6531.922047547547u,0 6531.923047547547u,1.5 6532.899587587588u,1.5 6532.900587587588u,0 6533.8771276276275u,0 6533.878127627628u,1.5 6534.854667667668u,1.5 6534.855667667668u,0 6535.832207707707u,0 6535.8332077077075u,1.5 6536.809747747748u,1.5 6536.810747747748u,0 6537.787287787788u,0 6537.788287787788u,1.5 6538.7648278278275u,1.5 6538.765827827828u,0 6539.742367867868u,0 6539.743367867868u,1.5 6545.607608108108u,1.5 6545.6086081081085u,0 6546.585148148148u,0 6546.586148148148u,1.5 6547.562688188188u,1.5 6547.563688188188u,0 6548.5402282282275u,0 6548.541228228228u,1.5 6550.495308308308u,1.5 6550.4963083083085u,0 6552.450388388388u,0 6552.451388388388u,1.5 6553.4279284284285u,1.5 6553.428928428429u,0 6554.405468468469u,0 6554.406468468469u,1.5 6555.383008508508u,1.5 6555.3840085085085u,0 6556.360548548548u,0 6556.361548548548u,1.5 6558.3156286286285u,1.5 6558.316628628629u,0 6560.270708708708u,0 6560.2717087087085u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6567.113488988989u,0 6567.114488988989u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.9787292292285u,0 6572.979729229229u,1.5 6573.95626926927u,1.5 6573.95726926927u,0 6575.911349349349u,0 6575.912349349349u,1.5 6577.866429429429u,1.5 6577.86742942943u,0 6578.84396946947u,0 6578.84496946947u,1.5 6579.821509509509u,1.5 6579.8225095095095u,0 6584.709209709709u,0 6584.7102097097095u,1.5 6588.61936986987u,1.5 6588.62036986987u,0 6592.5295300300295u,0 6592.53053003003u,1.5 6598.394770270271u,1.5 6598.395770270271u,0 6599.37231031031u,0 6599.37331031031u,1.5 6601.32739039039u,1.5 6601.32839039039u,0 6602.30493043043u,0 6602.305930430431u,1.5 6603.282470470471u,1.5 6603.283470470471u,0 6606.215090590591u,0 6606.216090590591u,1.5 6608.170170670671u,1.5 6608.171170670671u,0 6609.14771071071u,0 6609.1487107107105u,1.5 6614.03541091091u,1.5 6614.0364109109105u,0 6615.990490990991u,0 6615.991490990991u,1.5 6616.9680310310305u,1.5 6616.969031031031u,0 6619.900651151151u,0 6619.901651151151u,1.5 6620.878191191191u,1.5 6620.879191191191u,0 6622.833271271272u,0 6622.834271271272u,1.5 6623.810811311311u,1.5 6623.811811311311u,0 6624.788351351351u,0 6624.789351351351u,1.5 6629.676051551551u,1.5 6629.677051551551u,0 6630.653591591592u,0 6630.654591591592u,1.5 6633.586211711711u,1.5 6633.5872117117115u,0 6634.563751751752u,0 6634.564751751752u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6640.428991991992u,1.5 6640.429991991992u,0 6642.384072072072u,0 6642.385072072072u,1.5 6643.361612112112u,1.5 6643.362612112112u,0 6645.316692192192u,0 6645.317692192192u,1.5 6646.2942322322315u,1.5 6646.295232232232u,0 6650.204392392392u,0 6650.205392392392u,1.5 6652.159472472473u,1.5 6652.160472472473u,0 6654.114552552552u,0 6654.115552552552u,1.5 6655.092092592593u,1.5 6655.093092592593u,0 6656.069632632632u,0 6656.070632632633u,1.5 6657.047172672673u,1.5 6657.048172672673u,0 6658.024712712712u,0 6658.025712712712u,1.5 6659.002252752753u,1.5 6659.003252752753u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6666.822573073073u,1.5 6666.823573073073u,0 6667.800113113113u,0 6667.801113113113u,1.5 6668.777653153153u,1.5 6668.778653153153u,0 6671.710273273274u,0 6671.711273273274u,1.5 6672.687813313313u,1.5 6672.688813313313u,0 6674.642893393393u,0 6674.643893393393u,1.5 6676.597973473474u,1.5 6676.598973473474u,0 6677.575513513513u,0 6677.576513513513u,1.5 6678.553053553553u,1.5 6678.554053553553u,0 6679.530593593594u,0 6679.531593593594u,1.5 6680.508133633633u,1.5 6680.509133633634u,0 6684.418293793794u,0 6684.419293793794u,1.5 6685.395833833833u,1.5 6685.396833833834u,0 6687.350913913913u,0 6687.351913913913u,1.5 6689.305993993994u,1.5 6689.306993993994u,0 6690.283534034033u,0 6690.284534034034u,1.5 6692.238614114114u,1.5 6692.239614114114u,0 6697.126314314314u,0 6697.127314314314u,1.5 6702.991554554554u,1.5 6702.992554554554u,0 6707.879254754755u,0 6707.880254754755u,1.5 6710.811874874875u,1.5 6710.812874874875u,0 6711.789414914914u,0 6711.790414914914u,1.5 6712.766954954955u,1.5 6712.767954954955u,0 6713.744494994995u,0 6713.745494994995u,1.5 6714.722035035034u,1.5 6714.723035035035u,0 6715.699575075075u,0 6715.700575075075u,1.5 6717.654655155155u,1.5 6717.655655155155u,0 6719.609735235234u,0 6719.610735235235u,1.5 6720.587275275276u,1.5 6720.588275275276u,0 6724.497435435435u,0 6724.498435435436u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6729.385135635635u,0 6729.386135635636u,1.5 6730.362675675676u,1.5 6730.363675675676u,0 6731.340215715715u,0 6731.341215715715u,1.5 6734.272835835835u,1.5 6734.273835835836u,0 6735.250375875876u,0 6735.251375875876u,1.5 6736.227915915916u,1.5 6736.228915915916u,0 6739.160536036035u,0 6739.161536036036u,1.5 6740.138076076076u,1.5 6740.139076076076u,0 6741.115616116116u,0 6741.116616116116u,1.5 6742.093156156156u,1.5 6742.094156156156u,0 6743.070696196196u,0 6743.071696196196u,1.5 6745.025776276277u,1.5 6745.026776276277u,0 6746.980856356356u,0 6746.981856356356u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5 6755.778716716716u,1.5 6755.779716716716u,0 6756.7562567567575u,0 6756.757256756758u,1.5 6759.688876876877u,1.5 6759.689876876877u,0 6762.621496996997u,0 6762.622496996997u,1.5 6766.5316571571575u,1.5 6766.532657157158u,0 6770.441817317317u,0 6770.442817317317u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6776.3070575575575u,1.5 6776.308057557558u,0 6780.217217717717u,0 6780.218217717717u,1.5 6784.127377877878u,1.5 6784.128377877878u,0 6785.104917917918u,0 6785.105917917918u,1.5 6788.037538038037u,1.5 6788.038538038038u,0 6792.925238238237u,0 6792.926238238238u,1.5 6798.790478478479u,1.5 6798.791478478479u,0 6799.768018518518u,0 6799.769018518518u,1.5 6800.7455585585585u,1.5 6800.746558558559u,0 6802.700638638638u,0 6802.7016386386385u,1.5 6804.655718718718u,1.5 6804.656718718718u,0 6806.610798798799u,0 6806.611798798799u,1.5 6808.565878878879u,1.5 6808.566878878879u,0 6809.543418918919u,0 6809.544418918919u,1.5 6810.520958958959u,1.5 6810.52195895896u,0 6812.476039039038u,0 6812.477039039039u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6816.386199199199u,0 6816.387199199199u,1.5 6819.318819319319u,1.5 6819.319819319319u,0 6820.2963593593595u,0 6820.29735935936u,1.5 6821.273899399399u,1.5 6821.274899399399u,0 6823.22897947948u,0 6823.22997947948u,1.5 6825.1840595595595u,1.5 6825.18505955956u,0 6826.1615995996u,0 6826.1625995996u,1.5 6827.139139639639u,1.5 6827.1401396396395u,0 6828.11667967968u,0 6828.11767967968u,1.5 6831.0492997998u,1.5 6831.0502997998u,0 6832.026839839839u,0 6832.0278398398395u,1.5 6833.00437987988u,1.5 6833.00537987988u,0 6837.89208008008u,0 6837.89308008008u,1.5 6843.75732032032u,1.5 6843.75832032032u,0 6844.7348603603605u,0 6844.735860360361u,1.5 6845.7124004004u,1.5 6845.7134004004u,0 6846.68994044044u,0 6846.6909404404405u,1.5 6847.667480480481u,1.5 6847.668480480481u,0 6850.600100600601u,0 6850.601100600601u,1.5 6854.510260760761u,1.5 6854.511260760762u,0 6855.487800800801u,0 6855.488800800801u,1.5 6856.46534084084u,1.5 6856.4663408408405u,0 6857.442880880881u,0 6857.443880880881u,1.5 6859.397960960961u,1.5 6859.398960960962u,0 6864.285661161161u,0 6864.286661161162u,1.5 6865.263201201201u,1.5 6865.264201201201u,0 6866.24074124124u,0 6866.241741241241u,1.5 6872.105981481482u,1.5 6872.106981481482u,0 6873.083521521521u,0 6873.084521521521u,1.5 6874.0610615615615u,1.5 6874.062061561562u,0 6877.971221721721u,0 6877.972221721721u,1.5 6878.948761761762u,1.5 6878.949761761763u,0 6879.926301801802u,0 6879.927301801802u,1.5 6883.836461961962u,1.5 6883.837461961963u,0 6884.814002002002u,0 6884.815002002002u,1.5 6886.769082082082u,1.5 6886.770082082082u,0 6889.701702202202u,0 6889.702702202202u,1.5 6890.679242242241u,1.5 6890.680242242242u,0 6891.656782282283u,0 6891.657782282283u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5 6902.409722722722u,1.5 6902.410722722722u,0 6903.387262762763u,0 6903.388262762764u,1.5 6904.364802802803u,1.5 6904.365802802803u,0 6911.207583083083u,0 6911.208583083083u,1.5 6912.185123123123u,1.5 6912.186123123123u,0 6913.162663163163u,0 6913.163663163164u,1.5 6915.117743243242u,1.5 6915.1187432432425u,0 6916.095283283284u,0 6916.096283283284u,1.5 6918.050363363363u,1.5 6918.051363363364u,0 6919.027903403403u,0 6919.028903403403u,1.5 6921.960523523523u,1.5 6921.961523523523u,0 6924.893143643643u,0 6924.8941436436435u,1.5 6925.870683683684u,1.5 6925.871683683684u,0 6929.780843843843u,0 6929.7818438438435u,1.5 6930.758383883884u,1.5 6930.759383883884u,0 6935.646084084084u,0 6935.647084084084u,1.5 6937.601164164164u,1.5 6937.602164164165u,0 6938.578704204204u,0 6938.579704204204u,1.5 6943.466404404404u,1.5 6943.467404404404u,0 6945.421484484485u,0 6945.422484484485u,1.5 6946.399024524524u,1.5 6946.400024524524u,0 6947.376564564564u,0 6947.377564564565u,1.5 6949.331644644644u,1.5 6949.3326446446445u,0 6952.264264764765u,0 6952.265264764766u,1.5 6953.241804804805u,1.5 6953.242804804805u,0 6956.174424924925u,0 6956.175424924925u,1.5 6959.107045045044u,1.5 6959.1080450450445u,0 6963.994745245244u,0 6963.9957452452445u,1.5 6964.972285285286u,1.5 6964.973285285286u,0 6965.949825325325u,0 6965.950825325325u,1.5 6966.927365365365u,1.5 6966.928365365366u,0 6968.882445445445u,0 6968.883445445445u,1.5 6971.815065565565u,1.5 6971.816065565566u,0 6972.792605605606u,0 6972.793605605606u,1.5 6973.770145645645u,1.5 6973.771145645645u,0 6974.747685685686u,0 6974.748685685686u,1.5 6975.725225725725u,1.5 6975.726225725725u,0 6976.702765765766u,0 6976.703765765767u,1.5 6980.612925925926u,1.5 6980.613925925926u,0 6981.590465965966u,0 6981.591465965967u,1.5 6986.478166166166u,1.5 6986.479166166167u,0 6989.410786286287u,0 6989.411786286287u,1.5 6990.388326326326u,1.5 6990.389326326326u,0 6991.365866366366u,0 6991.366866366367u,1.5 6992.343406406406u,1.5 6992.344406406406u,0 6993.320946446446u,0 6993.321946446446u,1.5 6996.253566566566u,1.5 6996.254566566567u,0 6997.231106606607u,0 6997.232106606607u,1.5
vb22 b22 0 pwl 0,0  17.59522072072072u,0 17.59622072072072u,1.5 18.572760760760765u,1.5 18.573760760760763u,0 21.50538088088088u,0 21.50638088088088u,1.5 22.482920920920925u,1.5 22.483920920920923u,0 27.370621121121122u,0 27.37162112112112u,1.5 28.348161161161162u,1.5 28.34916116116116u,0 29.325701201201202u,0 29.3267012012012u,1.5 30.303241241241246u,1.5 30.304241241241243u,0 32.25832132132132u,0 32.25932132132132u,1.5 37.146021521521526u,1.5 37.14702152152153u,0 38.12356156156156u,0 38.12456156156156u,1.5 40.07864164164164u,1.5 40.07964164164164u,0 41.05618168168168u,0 41.05718168168168u,1.5 61.58452252252251u,1.5 61.58552252252252u,0 62.56206256256256u,0 62.563062562562564u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 64.51714264264264u,0 64.51814264264264u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 67.44976276276276u,1.5 67.45076276276276u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 70.38238288288288u,0 70.38338288288288u,1.5 71.35992292292292u,1.5 71.36092292292292u,0 81.13532332332332u,0 81.13632332332332u,1.5 82.11286336336336u,1.5 82.11386336336336u,0 85.04548348348348u,0 85.04648348348348u,1.5 86.02302352352352u,1.5 86.02402352352352u,0 88.95564364364364u,0 88.95664364364364u,1.5 89.9331836836837u,1.5 89.9341836836837u,0 90.91072372372372u,0 90.91172372372372u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 120.23692492492492u,0 120.23792492492493u,1.5 121.21446496496498u,1.5 121.21546496496498u,0 122.19200500500502u,0 122.19300500500502u,1.5 124.14708508508508u,1.5 124.14808508508509u,0 125.12462512512512u,0 125.12562512512513u,1.5 134.90002552552554u,1.5 134.9010255255255u,0 135.8775655655656u,0 135.87856556556557u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 148.58558608608612u,0 148.5865860860861u,1.5 149.56312612612612u,1.5 149.5641261261261u,0 150.54066616616618u,0 150.54166616616615u,1.5 151.51820620620623u,1.5 151.5192062062062u,0 152.49574624624626u,0 152.49674624624623u,1.5 163.2486866866867u,1.5 163.2496866866867u,0 174.00162712712714u,0 174.0026271271271u,1.5 177.9117872872873u,1.5 177.91278728728727u,0 178.88932732732735u,0 178.89032732732733u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 194.529967967968u,0 194.53096796796797u,1.5 195.50750800800802u,1.5 195.508508008008u,0 197.4625880880881u,0 197.46358808808807u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 217.0133888888889u,0 217.01438888888887u,1.5 217.99092892892892u,1.5 217.9919289289289u,0 218.96846896896898u,0 218.96946896896895u,1.5 221.90108908908908u,1.5 221.90208908908906u,0 222.87862912912914u,0 222.8796291291291u,1.5 225.81124924924927u,1.5 225.81224924924925u,0 226.7887892892893u,0 226.78978928928927u,1.5 228.74386936936938u,1.5 228.74486936936935u,0 239.4968098098098u,0 239.49780980980978u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 259.04761061061066u,0 259.04861061061064u,1.5 260.02515065065063u,1.5 260.0261506506506u,0 261.98023073073074u,0 261.9812307307307u,1.5 262.95777077077076u,1.5 262.95877077077074u,0 263.93531081081085u,0 263.9363108108108u,1.5 264.9128508508509u,1.5 264.91385085085085u,0 265.8903908908909u,0 265.8913908908909u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 280.5534914914915u,0 280.5544914914915u,1.5 281.53103153153154u,1.5 281.5320315315315u,0 282.50857157157157u,0 282.50957157157154u,1.5 283.48611161161165u,1.5 283.4871116116116u,0 284.4636516516517u,0 284.46465165165165u,1.5 291.3064319319319u,1.5 291.3074319319319u,0 292.28397197197194u,0 292.2849719719719u,1.5 294.23905205205205u,1.5 294.240052052052u,0 302.0593723723724u,0 302.0603723723724u,1.5 303.03691241241245u,1.5 303.0379124124124u,0 304.9919924924925u,0 304.9929924924925u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 316.722472972973u,0 316.72347297297296u,1.5 317.700013013013u,1.5 317.701013013013u,0 325.5203333333333u,0 325.5213333333333u,1.5 326.4978733733734u,1.5 326.4988733733734u,0 327.47541341341343u,0 327.4764134134134u,1.5 329.4304934934935u,1.5 329.43149349349346u,0 330.4080335335335u,0 330.4090335335335u,1.5 334.31819369369373u,1.5 334.3191936936937u,0 335.2957337337337u,0 335.2967337337337u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 348.9812942942943u,0 348.98229429429426u,1.5 349.9588343343343u,1.5 349.9598343343343u,0 350.9363743743744u,0 350.9373743743744u,1.5 351.9139144144144u,1.5 351.9149144144144u,0 352.8914544544545u,0 352.8924544544545u,1.5 353.8689944944945u,1.5 353.86999449449445u,0 354.8465345345345u,0 354.8475345345345u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 377.3299554554555u,0 377.33095545545547u,1.5 378.3074954954955u,1.5 378.3084954954955u,0 379.28503553553554u,0 379.2860355355355u,1.5 391.99305605605605u,1.5 391.994056056056u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 406.65615665665666u,0 406.65715665665664u,1.5 407.6336966966967u,1.5 407.63469669669666u,0 409.5887767767768u,0 409.5897767767768u,1.5 410.5663168168168u,1.5 410.5673168168168u,0 413.49893693693696u,0 413.49993693693693u,1.5 416.43155705705703u,1.5 416.432557057057u,0 417.40909709709706u,0 417.41009709709704u,1.5 434.0272777777778u,1.5 434.02827777777776u,0 435.98235785785783u,0 435.9833578578578u,1.5 436.9598978978979u,1.5 436.9608978978979u,0 442.82513813813813u,0 442.8261381381381u,1.5 443.80267817817816u,1.5 443.80367817817813u,0 447.7128383383383u,0 447.7138383383383u,1.5 448.69037837837834u,1.5 448.6913783783783u,0 462.37593893893893u,0 462.3769389389389u,1.5 463.353478978979u,1.5 463.354478978979u,0 467.2636391391391u,0 467.2646391391391u,1.5 468.2411791791792u,1.5 468.2421791791792u,0 470.19625925925925u,0 470.1972592592592u,1.5 472.15133933933936u,1.5 472.15233933933933u,0 473.1288793793794u,0 473.12987937937936u,1.5 474.1064194194194u,1.5 474.1074194194194u,0 475.08395945945944u,0 475.0849594594594u,1.5 478.0165795795796u,1.5 478.0175795795796u,0 478.9941196196196u,0 478.9951196196196u,1.5 481.92673973973973u,1.5 481.9277397397397u,0 482.9042797797798u,0 482.9052797797798u,1.5 484.8593598598599u,1.5 484.8603598598599u,0 485.8368998998999u,0 485.83789989989987u,1.5 489.7470600600601u,1.5 489.7480600600601u,0 490.72460010010013u,0 490.7256001001001u,1.5 512.2304809809809u,1.5 512.2314809809809u,0 513.2080210210211u,0 513.209021021021u,1.5 514.1855610610611u,1.5 514.1865610610611u,0 515.1631011011011u,0 515.1641011011011u,1.5 516.1406411411411u,1.5 516.1416411411411u,0 517.1181811811812u,0 517.1191811811811u,1.5 518.0957212212213u,1.5 518.0967212212213u,0 519.0732612612613u,0 519.0742612612613u,1.5 520.0508013013012u,1.5 520.0518013013012u,0 521.0283413413413u,0 521.0293413413413u,1.5 525.9160415415415u,1.5 525.9170415415415u,0 526.8935815815815u,0 526.8945815815815u,1.5 527.8711216216217u,1.5 527.8721216216217u,0 529.8262017017017u,0 529.8272017017017u,1.5 531.7812817817818u,1.5 531.7822817817818u,0 534.7139019019019u,0 534.7149019019018u,1.5 535.6914419419419u,1.5 535.6924419419419u,0 537.646522022022u,0 537.647522022022u,1.5 538.6240620620621u,1.5 538.625062062062u,0 560.1299429429429u,0 560.1309429429429u,1.5 562.085023023023u,1.5 562.086023023023u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 567.9502632632633u,1.5 567.9512632632633u,0 568.9278033033033u,0 568.9288033033033u,1.5 587.501064064064u,1.5 587.502064064064u,0 588.4786041041041u,0 588.479604104104u,1.5 589.4561441441441u,1.5 589.4571441441441u,0 591.4112242242243u,0 591.4122242242242u,1.5 592.3887642642643u,1.5 592.3897642642643u,0 605.0967847847849u,0 605.0977847847848u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 608.0294049049048u,0 608.0304049049048u,1.5 619.7598853853854u,1.5 619.7608853853853u,0 620.7374254254254u,0 620.7384254254254u,1.5 621.7149654654654u,1.5 621.7159654654654u,0 622.6925055055054u,0 622.6935055055054u,1.5 623.6700455455456u,1.5 623.6710455455456u,0 633.445445945946u,0 633.4464459459459u,1.5 634.422985985986u,1.5 634.423985985986u,0 635.400526026026u,0 635.401526026026u,1.5 636.378066066066u,1.5 636.379066066066u,0 637.355606106106u,0 637.356606106106u,1.5 646.1534664664664u,1.5 646.1544664664664u,0 647.1310065065064u,0 647.1320065065064u,1.5 650.0636266266266u,1.5 650.0646266266266u,0 661.7941071071072u,0 661.7951071071071u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 665.7042672672673u,0 665.7052672672672u,1.5 673.5245875875876u,1.5 673.5255875875876u,0 674.5021276276276u,0 674.5031276276276u,1.5 675.4796676676676u,1.5 675.4806676676676u,0 678.4122877877878u,0 678.4132877877878u,1.5 679.3898278278278u,1.5 679.3908278278278u,0 684.277528028028u,0 684.278528028028u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 696.9855485485485u,1.5 696.9865485485485u,0 697.9630885885886u,0 697.9640885885885u,1.5 698.9406286286286u,1.5 698.9416286286286u,0 704.8058688688689u,0 704.8068688688688u,1.5 705.783408908909u,1.5 705.784408908909u,0 708.716029029029u,0 708.7170290290289u,1.5 718.4914294294294u,1.5 718.4924294294294u,0 719.4689694694696u,0 719.4699694694696u,1.5 720.4465095095095u,1.5 720.4475095095095u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 730.22190990991u,0 730.22290990991u,1.5 739.0197702702703u,1.5 739.0207702702703u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 758.5705710710711u,1.5 758.571571071071u,0 759.5481111111111u,0 759.5491111111111u,1.5 761.5031911911911u,1.5 761.5041911911911u,0 763.4582712712713u,0 763.4592712712713u,1.5 764.4358113113113u,1.5 764.4368113113113u,0 770.3010515515515u,0 770.3020515515515u,1.5 780.076451951952u,1.5 780.077451951952u,0 781.053991991992u,0 781.054991991992u,1.5 783.0090720720721u,1.5 783.010072072072u,0 791.8069324324325u,0 791.8079324324325u,1.5 801.5823328328329u,1.5 801.5833328328329u,0 802.5598728728729u,0 802.5608728728729u,1.5 803.5374129129129u,1.5 803.5384129129129u,0 804.514952952953u,0 804.515952952953u,1.5 805.492492992993u,1.5 805.493492992993u,0 813.3128133133133u,0 813.3138133133133u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 816.2454334334335u,0 816.2464334334335u,1.5 817.2229734734735u,1.5 817.2239734734735u,0 818.2005135135136u,0 818.2015135135135u,1.5 825.0432937937937u,1.5 825.0442937937937u,0 826.0208338338339u,0 826.0218338338339u,1.5 826.9983738738739u,1.5 826.9993738738739u,0 834.8186941941941u,0 834.8196941941941u,1.5 835.7962342342342u,1.5 835.7972342342342u,0 836.7737742742743u,0 836.7747742742743u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 849.4817947947948u,1.5 849.4827947947948u,0 850.4593348348349u,0 850.4603348348348u,1.5 851.4368748748749u,1.5 851.4378748748749u,0 853.3919549549549u,0 853.3929549549549u,1.5 854.3694949949951u,1.5 854.370494994995u,0 861.2122752752753u,0 861.2132752752752u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 866.0999754754755u,0 866.1009754754755u,1.5 874.8978358358358u,1.5 874.8988358358358u,0 875.8753758758759u,0 875.8763758758759u,1.5 877.8304559559559u,1.5 877.8314559559559u,0 878.8079959959961u,0 878.808995995996u,1.5 879.7855360360361u,1.5 879.7865360360361u,0 895.4261766766766u,0 895.4271766766766u,1.5 905.2015770770771u,1.5 905.2025770770771u,0 906.1791171171171u,0 906.1801171171171u,1.5 910.0892772772772u,1.5 910.0902772772772u,0 911.0668173173173u,0 911.0678173173172u,1.5 912.0443573573574u,1.5 912.0453573573574u,0 913.9994374374375u,0 914.0004374374374u,1.5 914.9769774774775u,1.5 914.9779774774775u,0 918.8871376376377u,0 918.8881376376377u,1.5 919.8646776776777u,1.5 919.8656776776777u,0 929.6400780780781u,0 929.6410780780781u,1.5 930.6176181181181u,1.5 930.6186181181181u,0 934.5277782782782u,0 934.5287782782782u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 936.4828583583584u,0 936.4838583583584u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 940.3930185185185u,0 940.3940185185185u,1.5 961.8988993993994u,1.5 961.8998993993994u,0 962.8764394394394u,0 962.8774394394394u,1.5 964.8315195195195u,1.5 964.8325195195195u,0 965.8090595595596u,0 965.8100595595596u,1.5 968.7416796796797u,1.5 968.7426796796797u,0 970.6967597597597u,0 970.6977597597597u,1.5 972.6518398398398u,1.5 972.6528398398398u,0 973.6293798798798u,0 973.6303798798798u,1.5 974.60691991992u,1.5 974.6079199199199u,0 975.58445995996u,0 975.58545995996u,1.5 976.562u,1.5 976.563u,0 977.5395400400402u,0 977.5405400400401u,1.5 978.5170800800801u,1.5 978.51808008008u,0 982.4272402402403u,0 982.4282402402403u,1.5 983.4047802802802u,1.5 983.4057802802802u,0 984.3823203203203u,0 984.3833203203203u,1.5 985.3598603603602u,1.5 985.3608603603602u,0 988.2924804804804u,0 988.2934804804804u,1.5 989.2700205205206u,1.5 989.2710205205206u,0 999.045420920921u,0 999.0464209209209u,1.5 1000.0229609609609u,1.5 1000.0239609609608u,0 1001.000501001001u,0 1001.001501001001u,1.5 1001.9780410410411u,1.5 1001.9790410410411u,0 1011.7534414414415u,0 1011.7544414414415u,1.5 1012.7309814814814u,1.5 1012.7319814814814u,0 1013.7085215215216u,0 1013.7095215215215u,1.5 1014.6860615615615u,1.5 1014.6870615615614u,0 1021.5288418418419u,0 1021.5298418418419u,1.5 1022.5063818818818u,1.5 1022.5073818818818u,0 1023.4839219219219u,0 1023.4849219219219u,1.5 1025.4390020020019u,1.5 1025.440002002002u,0 1026.416542042042u,0 1026.4175420420422u,1.5 1027.394082082082u,1.5 1027.3950820820821u,0 1028.371622122122u,0 1028.3726221221223u,1.5 1029.349162162162u,1.5 1029.3501621621622u,0 1030.3267022022021u,0 1030.3277022022023u,1.5 1031.3042422422423u,1.5 1031.3052422422425u,0 1032.2817822822822u,0 1032.2827822822824u,1.5 1034.2368623623622u,1.5 1034.2378623623624u,0 1035.2144024024024u,0 1035.2154024024026u,1.5 1038.1470225225225u,1.5 1038.1480225225228u,0 1039.1245625625625u,0 1039.1255625625627u,1.5 1063.5630635635634u,1.5 1063.5640635635636u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1085.0689444444445u,0 1085.0699444444447u,1.5 1086.0464844844844u,1.5 1086.0474844844846u,0 1087.0240245245245u,0 1087.0250245245247u,1.5 1088.9791046046046u,1.5 1088.9801046046048u,0 1089.9566446446445u,0 1089.9576446446447u,1.5 1091.9117247247245u,1.5 1091.9127247247247u,0 1092.8892647647647u,0 1092.8902647647649u,1.5 1094.8443448448447u,1.5 1094.845344844845u,0 1095.8218848848846u,0 1095.8228848848848u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1120.2603858858856u,0 1120.2613858858858u,1.5 1121.2379259259258u,1.5 1121.238925925926u,0 1122.215465965966u,0 1122.216465965966u,1.5 1123.1930060060058u,1.5 1123.194006006006u,0 1124.170546046046u,0 1124.1715460460462u,1.5 1126.125626126126u,1.5 1126.1266261261262u,0 1127.1031661661661u,0 1127.1041661661664u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1137.8561066066065u,1.5 1137.8571066066067u,0 1148.609047047047u,0 1148.6100470470471u,1.5 1149.5865870870869u,1.5 1149.587587087087u,0 1150.564127127127u,0 1150.5651271271272u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1174.0250880880878u,0 1174.026088088088u,1.5 1175.9801681681681u,1.5 1175.9811681681683u,0 1176.957708208208u,0 1176.9587082082082u,1.5 1182.8229484484484u,1.5 1182.8239484484486u,0 1183.8004884884883u,0 1183.8014884884885u,1.5 1184.7780285285285u,1.5 1184.7790285285287u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1186.7331086086085u,1.5 1186.7341086086087u,0 1195.5309689689689u,0 1195.531968968969u,1.5 1196.5085090090088u,1.5 1196.509509009009u,0 1197.486049049049u,0 1197.4870490490491u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1214.1042297297297u,0 1214.10522972973u,1.5 1215.0817697697696u,1.5 1215.0827697697698u,0 1217.0368498498497u,0 1217.0378498498499u,1.5 1218.0143898898898u,1.5 1218.01538988989u,0 1218.9919299299297u,0 1218.99292992993u,1.5 1227.7897902902903u,1.5 1227.7907902902905u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1239.5202707707706u,0 1239.5212707707708u,1.5 1241.4753508508506u,1.5 1241.4763508508508u,0 1242.4528908908908u,0 1242.453890890891u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1259.0710715715716u,0 1259.0720715715718u,1.5 1261.0261516516516u,1.5 1261.0271516516518u,0 1262.0036916916918u,0 1262.004691691692u,1.5 1264.9363118118117u,1.5 1264.937311811812u,0 1265.9138518518516u,0 1265.9148518518518u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1269.8240120120117u,0 1269.825012012012u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1282.5320325325324u,0 1282.5330325325326u,1.5 1289.3748128128127u,1.5 1289.375812812813u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1295.2400530530529u,1.5 1295.241053053053u,0 1299.150213213213u,0 1299.1512132132132u,1.5 1300.127753253253u,1.5 1300.1287532532533u,0 1301.1052932932932u,0 1301.1062932932934u,1.5 1302.0828333333332u,1.5 1302.0838333333334u,0 1303.0603733733733u,0 1303.0613733733735u,1.5 1305.0154534534533u,1.5 1305.0164534534536u,0 1305.9929934934935u,0 1305.9939934934937u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1324.566254254254u,0 1324.5672542542543u,1.5 1325.5437942942942u,1.5 1325.5447942942944u,0 1326.5213343343341u,0 1326.5223343343343u,1.5 1336.2967347347346u,1.5 1336.2977347347348u,0 1337.2742747747748u,0 1337.275274774775u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1340.2068948948947u,0 1340.207894894895u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1350.9598353353351u,0 1350.9608353353353u,1.5 1352.9149154154154u,1.5 1352.9159154154156u,0 1353.8924554554553u,0 1353.8934554554555u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1363.6678558558558u,1.5 1363.668855855856u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1365.6229359359356u,1.5 1365.6239359359358u,0 1378.3309564564563u,0 1378.3319564564565u,1.5 1380.2860365365364u,1.5 1380.2870365365366u,0 1381.2635765765765u,0 1381.2645765765767u,1.5 1391.0389769769768u,1.5 1391.039976976977u,0 1392.016517017017u,0 1392.017517017017u,1.5 1392.9940570570568u,1.5 1392.995057057057u,0 1393.971597097097u,0 1393.9725970970972u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1395.926677177177u,0 1395.9276771771772u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1408.6346976976977u,0 1408.6356976976979u,1.5 1409.6122377377376u,1.5 1409.6132377377378u,0 1412.5448578578578u,0 1412.545857857858u,1.5 1413.522397897898u,1.5 1413.5233978978981u,0 1415.4774779779777u,0 1415.478477977978u,1.5 1416.4550180180179u,1.5 1416.456018018018u,0 1417.4325580580578u,0 1417.433558058058u,1.5 1418.410098098098u,1.5 1418.4110980980981u,0 1419.3876381381378u,0 1419.388638138138u,1.5 1436.9833588588588u,1.5 1436.984358858859u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1440.8935190190189u,1.5 1440.894519019019u,0 1441.8710590590588u,0 1441.872059059059u,1.5 1442.848599099099u,1.5 1442.8495990990991u,0 1448.7138393393393u,0 1448.7148393393395u,1.5 1449.6913793793792u,1.5 1449.6923793793794u,0 1463.37693993994u,0 1463.3779399399402u,1.5 1464.35447997998u,1.5 1464.3554799799801u,0 1466.3095600600598u,0 1466.31056006006u,1.5 1467.2871001001u,1.5 1467.2881001001u,0 1468.26464014014u,0 1468.2656401401402u,1.5 1469.24218018018u,1.5 1469.2431801801802u,0 1473.1523403403403u,0 1473.1533403403405u,1.5 1474.1298803803802u,1.5 1474.1308803803804u,0 1476.0849604604603u,0 1476.0859604604605u,1.5 1478.0400405405405u,1.5 1478.0410405405407u,0 1479.0175805805804u,0 1479.0185805805806u,1.5 1482.9277407407408u,1.5 1482.928740740741u,0 1483.9052807807807u,0 1483.906280780781u,1.5 1486.8379009009009u,1.5 1486.838900900901u,0 1487.815440940941u,0 1487.8164409409412u,1.5 1494.658221221221u,1.5 1494.6592212212213u,0 1495.635761261261u,0 1495.6367612612612u,1.5 1497.5908413413413u,1.5 1497.5918413413415u,0 1498.5683813813812u,0 1498.5693813813814u,1.5 1499.5459214214213u,1.5 1499.5469214214215u,0 1500.5234614614612u,0 1500.5244614614614u,1.5 1506.3887017017016u,1.5 1506.3897017017018u,0 1507.3662417417418u,0 1507.367241741742u,1.5 1512.253941941942u,1.5 1512.2549419419422u,0 1513.231481981982u,0 1513.2324819819821u,1.5 1514.209022022022u,1.5 1514.2100220220223u,0 1515.186562062062u,0 1515.1875620620622u,1.5 1521.0518023023021u,1.5 1521.0528023023023u,0 1522.0293423423423u,0 1522.0303423423425u,1.5 1525.9395025025024u,1.5 1525.9405025025026u,0 1528.8721226226226u,0 1528.8731226226228u,1.5 1529.8496626626625u,1.5 1529.8506626626627u,0 1530.8272027027026u,0 1530.8282027027028u,1.5 1531.8047427427427u,1.5 1531.805742742743u,0 1534.7373628628627u,0 1534.738362862863u,1.5 1535.7149029029028u,1.5 1535.715902902903u,0 1537.669982982983u,0 1537.670982982983u,1.5 1538.647523023023u,1.5 1538.6485230230232u,0 1540.6026031031029u,0 1540.603603103103u,1.5 1541.580143143143u,1.5 1541.5811431431432u,0 1561.130943943944u,0 1561.1319439439442u,1.5 1562.108483983984u,1.5 1562.109483983984u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1566.018644144144u,1.5 1566.0196441441442u,0 1566.996184184184u,0 1566.997184184184u,1.5 1583.614364864865u,1.5 1583.6153648648651u,0 1584.5919049049048u,0 1584.592904904905u,1.5 1587.524525025025u,1.5 1587.5255250250252u,0 1589.479605105105u,0 1589.4806051051053u,1.5 1590.457145145145u,1.5 1590.4581451451452u,0 1601.2100855855854u,0 1601.2110855855856u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1608.052865865866u,0 1608.053865865866u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1619.7833463463462u,1.5 1619.7843463463464u,0 1620.7608863863861u,0 1620.7618863863863u,1.5 1621.7384264264263u,1.5 1621.7394264264265u,0 1622.7159664664664u,0 1622.7169664664666u,1.5 1623.6935065065063u,1.5 1623.6945065065065u,0 1624.6710465465464u,0 1624.6720465465467u,1.5 1625.6485865865864u,1.5 1625.6495865865866u,0 1633.4689069069068u,0 1633.469906906907u,1.5 1634.446446946947u,1.5 1634.4474469469471u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1639.3341471471472u,1.5 1639.3351471471474u,0 1640.311687187187u,0 1640.3126871871873u,1.5 1649.1095475475474u,1.5 1649.1105475475476u,0 1651.0646276276275u,0 1651.0656276276277u,1.5 1652.0421676676676u,1.5 1652.0431676676678u,0 1658.884947947948u,0 1658.8859479479481u,1.5 1659.8624879879878u,1.5 1659.863487987988u,0 1663.7726481481482u,0 1663.7736481481484u,1.5 1674.5255885885883u,1.5 1674.5265885885885u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1686.256069069069u,1.5 1686.2570690690693u,0 1687.233609109109u,0 1687.2346091091092u,1.5 1696.0314694694694u,1.5 1696.0324694694696u,0 1697.9865495495494u,0 1697.9875495495496u,1.5 1698.9640895895895u,1.5 1698.9650895895898u,0 1706.7844099099098u,0 1706.78540990991u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1708.73948998999u,0 1708.7404899899902u,1.5 1711.67211011011u,1.5 1711.6731101101102u,0 1712.6496501501501u,0 1712.6506501501503u,1.5 1717.5373503503502u,1.5 1717.5383503503504u,0 1718.5148903903903u,0 1718.5158903903905u,1.5 1719.4924304304302u,1.5 1719.4934304304304u,0 1725.3576706706706u,0 1725.3586706706708u,1.5 1726.3352107107105u,1.5 1726.3362107107107u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1731.2229109109107u,1.5 1731.223910910911u,0 1732.2004509509509u,0 1732.201450950951u,1.5 1739.0432312312312u,1.5 1739.0442312312314u,0 1740.0207712712713u,0 1740.0217712712715u,1.5 1740.998311311311u,1.5 1740.9993113113112u,0 1741.9758513513511u,0 1741.9768513513513u,1.5 1742.9533913913913u,1.5 1742.9543913913915u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1760.549112112112u,1.5 1760.5501121121122u,0 1770.3245125125122u,0 1770.3255125125124u,1.5 1772.2795925925925u,1.5 1772.2805925925927u,0 1773.2571326326324u,0 1773.2581326326326u,1.5 1774.2346726726726u,1.5 1774.2356726726728u,0 1775.2122127127125u,0 1775.2132127127127u,1.5 1782.054992992993u,1.5 1782.0559929929932u,0 1791.8303933933933u,0 1791.8313933933935u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1800.6282537537536u,1.5 1800.6292537537538u,0 1801.6057937937937u,0 1801.606793793794u,1.5 1804.5384139139137u,1.5 1804.539413913914u,0 1811.3811941941942u,0 1811.3821941941944u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1814.3138143143142u,1.5 1814.3148143143144u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1823.1116746746745u,1.5 1823.1126746746747u,0 1824.0892147147147u,0 1824.0902147147149u,1.5 1826.0442947947947u,1.5 1826.045294794795u,0 1827.9993748748748u,0 1828.000374874875u,1.5 1828.976914914915u,1.5 1828.9779149149151u,0 1834.842155155155u,0 1834.8431551551553u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1851.4603358358356u,1.5 1851.4613358358358u,0 1861.235736236236u,0 1861.2367362362363u,1.5 1862.2132762762762u,1.5 1862.2142762762765u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1876.8763768768767u,1.5 1876.877376876877u,0 1877.853916916917u,0 1877.854916916917u,1.5 1878.8314569569568u,1.5 1878.832456956957u,0 1880.7865370370369u,0 1880.787537037037u,1.5 1881.764077077077u,1.5 1881.7650770770772u,0 1887.6293173173174u,0 1887.6303173173176u,1.5 1888.6068573573573u,1.5 1888.6078573573575u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1891.5394774774772u,1.5 1891.5404774774775u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1895.4496376376374u,0 1895.4506376376376u,1.5 1913.0453583583583u,1.5 1913.0463583583585u,0 1914.0228983983984u,0 1914.0238983983986u,1.5 1915.0004384384383u,1.5 1915.0014384384385u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1934.551239239239u,0 1934.5522392392393u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1939.4389394394395u,0 1939.4399394394397u,1.5 1960.94482032032u,1.5 1960.9458203203203u,0 1961.9223603603602u,0 1961.9233603603604u,1.5 1967.7876006006004u,1.5 1967.7886006006006u,0 1969.7426806806807u,0 1969.7436806806809u,1.5 1970.7202207207204u,1.5 1970.7212207207206u,0 1971.6977607607605u,0 1971.6987607607607u,1.5 1972.6753008008006u,1.5 1972.6763008008008u,0 1973.6528408408408u,0 1973.653840840841u,1.5 1974.630380880881u,1.5 1974.6313808808811u,0 1975.6079209209206u,0 1975.6089209209208u,1.5 1976.5854609609607u,1.5 1976.586460960961u,0 1978.540541041041u,0 1978.5415410410412u,1.5 1979.5180810810812u,1.5 1979.5190810810814u,0 1988.3159414414415u,0 1988.3169414414417u,1.5 1989.2934814814816u,1.5 1989.2944814814819u,0 1997.1138018018016u,0 1997.1148018018018u,1.5 1998.0913418418418u,1.5 1998.092341841842u,0 2002.979042042042u,0 2002.9800420420422u,1.5 2003.9565820820822u,1.5 2003.9575820820824u,0 2005.911662162162u,0 2005.9126621621622u,1.5 2006.8892022022021u,1.5 2006.8902022022023u,0 2017.6421426426425u,0 2017.6431426426427u,1.5 2018.6196826826827u,1.5 2018.6206826826829u,0 2020.5747627627625u,0 2020.5757627627627u,1.5 2021.5523028028026u,1.5 2021.5533028028028u,0 2024.4849229229226u,0 2024.4859229229228u,1.5 2025.4624629629627u,1.5 2025.463462962963u,0 2027.417543043043u,0 2027.4185430430432u,1.5 2030.350163163163u,1.5 2030.3511631631632u,0 2031.327703203203u,0 2031.3287032032033u,1.5 2032.3052432432432u,1.5 2032.3062432432434u,0 2033.2827832832834u,0 2033.2837832832836u,1.5 2038.1704834834836u,1.5 2038.1714834834838u,0 2039.1480235235233u,0 2039.1490235235235u,1.5 2058.698824324324u,1.5 2058.6998243243243u,0 2059.676364364364u,0 2059.677364364364u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2065.5416046046043u,0 2065.5426046046045u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2069.4517647647644u,1.5 2069.4527647647647u,0 2072.384384884885u,0 2072.3853848848853u,1.5 2073.3619249249246u,1.5 2073.3629249249248u,0 2088.025025525525u,0 2088.0260255255253u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2107.575826326326u,0 2107.576826326326u,1.5 2108.553366366366u,1.5 2108.554366366366u,0 2112.463526526526u,0 2112.4645265265262u,1.5 2113.4410665665664u,1.5 2113.4420665665666u,0 2122.2389269269265u,0 2122.2399269269267u,1.5 2123.216466966967u,1.5 2123.217466966967u,0 2124.194007007007u,0 2124.195007007007u,1.5 2125.171547047047u,1.5 2125.1725470470474u,0 2126.149087087087u,0 2126.1500870870873u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2147.654967967968u,0 2147.655967967968u,1.5 2148.632508008008u,1.5 2148.633508008008u,0 2149.610048048048u,0 2149.6110480480484u,1.5 2161.3405285285285u,1.5 2161.3415285285287u,0 2166.228228728729u,0 2166.229228728729u,1.5 2167.2057687687684u,1.5 2167.2067687687686u,0 2172.093468968969u,0 2172.094468968969u,1.5 2173.071009009009u,1.5 2173.072009009009u,0 2175.026089089089u,0 2175.0270890890893u,1.5 2177.9587092092092u,1.5 2177.9597092092094u,0 2178.936249249249u,0 2178.9372492492494u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2196.53196996997u,0 2196.53296996997u,1.5 2198.48705005005u,1.5 2198.4880500500503u,0 2199.46459009009u,0 2199.4655900900902u,1.5 2201.41967017017u,1.5 2201.42067017017u,0 2202.3972102102102u,0 2202.3982102102104u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2219.015390890891u,0 2219.016390890891u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2232.700951451451u,0 2232.7019514514514u,1.5 2233.6784914914915u,1.5 2233.6794914914917u,0 2240.5212717717714u,0 2240.5222717717716u,1.5 2241.4988118118117u,1.5 2241.499811811812u,0 2242.4763518518516u,0 2242.477351851852u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2258.1169924924925u,0 2258.1179924924927u,1.5 2259.0945325325324u,1.5 2259.0955325325326u,0 2261.0496126126122u,0 2261.0506126126124u,1.5 2262.0271526526526u,1.5 2262.028152652653u,0 2263.0046926926925u,0 2263.0056926926927u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2271.802553053053u,0 2271.8035530530533u,1.5 2272.780093093093u,1.5 2272.781093093093u,0 2281.577953453453u,0 2281.5789534534533u,1.5 2291.3533538538536u,1.5 2291.354353853854u,0 2292.330893893894u,0 2292.331893893894u,1.5 2294.285973973974u,1.5 2294.286973973974u,0 2304.0613743743743u,0 2304.0623743743745u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2317.746934934935u,0 2317.747934934935u,1.5 2318.724474974975u,1.5 2318.725474974975u,0 2326.5447952952954u,0 2326.5457952952956u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2348.050676176176u,0 2348.051676176176u,1.5 2349.028216216216u,1.5 2349.0292162162164u,0 2350.9832962962964u,0 2350.9842962962966u,1.5 2353.915916416416u,1.5 2353.9169164164164u,0 2354.893456456456u,0 2354.8944564564563u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2361.736236736737u,0 2361.737236736737u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2365.646396896897u,1.5 2365.647396896897u,0 2378.354417417417u,0 2378.3554174174174u,1.5 2379.331957457457u,1.5 2379.3329574574573u,0 2380.3094974974974u,0 2380.3104974974976u,1.5 2388.1298178178176u,1.5 2388.130817817818u,0 2389.1073578578576u,0 2389.1083578578578u,1.5 2393.0175180180177u,1.5 2393.018518018018u,0 2393.995058058058u,0 2393.996058058058u,1.5 2394.972598098098u,1.5 2394.973598098098u,0 2395.9501381381383u,0 2395.9511381381385u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2398.882758258258u,0 2398.8837582582582u,1.5 2399.8602982982984u,1.5 2399.8612982982986u,0 2408.6581586586585u,0 2408.6591586586587u,1.5 2409.6356986986984u,1.5 2409.6366986986986u,0 2413.5458588588585u,0 2413.5468588588587u,1.5 2430.1640395395393u,1.5 2430.1650395395395u,0 2431.1415795795797u,0 2431.14257957958u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.0068198198196u,0 2437.00781981982u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2463.400400900901u,0 2463.401400900901u,1.5 2465.355480980981u,1.5 2465.3564809809814u,0 2466.3330210210206u,0 2466.334021021021u,1.5 2467.310561061061u,1.5 2467.311561061061u,0 2469.2656411411413u,0 2469.2666411411415u,1.5 2470.243181181181u,1.5 2470.2441811811814u,0 2472.198261261261u,0 2472.199261261261u,1.5 2473.1758013013014u,1.5 2473.1768013013016u,0 2475.1308813813816u,0 2475.131881381382u,1.5 2476.108421421421u,1.5 2476.1094214214213u,0 2477.0859614614615u,0 2477.0869614614617u,1.5 2480.0185815815817u,1.5 2480.019581581582u,0 2480.996121621621u,0 2480.9971216216213u,1.5 2484.9062817817817u,1.5 2484.907281781782u,0 2485.8838218218216u,0 2485.884821821822u,1.5 2487.838901901902u,1.5 2487.839901901902u,0 2488.816441941942u,0 2488.817441941942u,1.5 2494.681682182182u,1.5 2494.6826821821824u,0 2495.659222222222u,0 2495.6602222222223u,1.5 2502.5020025025024u,1.5 2502.5030025025026u,0 2503.4795425425427u,0 2503.480542542543u,1.5 2504.4570825825826u,1.5 2504.458082582583u,0 2505.434622622622u,0 2505.4356226226223u,1.5 2507.3897027027024u,1.5 2507.3907027027026u,0 2508.3672427427427u,0 2508.368242742743u,1.5 2511.2998628628625u,1.5 2511.3008628628627u,0 2512.277402902903u,0 2512.278402902903u,1.5 2513.2549429429428u,1.5 2513.255942942943u,0 2514.232482982983u,0 2514.2334829829833u,1.5 2515.2100230230226u,1.5 2515.211023023023u,0 2516.187563063063u,0 2516.188563063063u,1.5 2522.0528033033033u,1.5 2522.0538033033035u,0 2523.0303433433432u,0 2523.0313433433435u,1.5 2524.0078833833836u,1.5 2524.008883383384u,0 2524.985423423423u,0 2524.9864234234233u,1.5 2526.9405035035034u,1.5 2526.9415035035036u,0 2527.9180435435437u,0 2527.919043543544u,1.5 2528.8955835835836u,1.5 2528.896583583584u,0 2530.8506636636635u,0 2530.8516636636637u,1.5 2531.8282037037034u,1.5 2531.8292037037036u,0 2532.8057437437437u,0 2532.806743743744u,1.5 2533.7832837837836u,1.5 2533.784283783784u,0 2535.7383638638635u,0 2535.7393638638637u,1.5 2536.715903903904u,1.5 2536.716903903904u,0 2540.626064064064u,0 2540.627064064064u,1.5 2541.603604104104u,1.5 2541.604604104104u,0 2563.109484984985u,0 2563.1104849849853u,1.5 2564.0870250250246u,1.5 2564.0880250250248u,0 2566.042105105105u,0 2566.043105105105u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2571.907345345345u,0 2571.9083453453454u,1.5 2579.7276656656654u,1.5 2579.7286656656656u,0 2580.7052057057053u,0 2580.7062057057055u,1.5 2581.6827457457457u,1.5 2581.683745745746u,0 2582.6602857857856u,0 2582.661285785786u,1.5 2588.5255260260255u,1.5 2588.5265260260257u,0 2590.480606106106u,0 2590.481606106106u,1.5 2591.458146146146u,1.5 2591.4591461461464u,0 2592.435686186186u,0 2592.4366861861863u,1.5 2593.413226226226u,1.5 2593.414226226226u,0 2601.2335465465467u,0 2601.234546546547u,1.5 2602.2110865865866u,1.5 2602.212086586587u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2607.0987867867866u,0 2607.099786786787u,1.5 2620.784347347347u,1.5 2620.7853473473474u,0 2623.7169674674674u,0 2623.7179674674676u,1.5 2624.6945075075073u,1.5 2624.6955075075075u,0 2625.6720475475477u,0 2625.673047547548u,1.5 2626.6495875875876u,1.5 2626.650587587588u,0 2636.424987987988u,0 2636.4259879879883u,1.5 2638.380068068068u,1.5 2638.381068068068u,0 2639.357608108108u,0 2639.358608108108u,1.5 2648.1554684684684u,1.5 2648.1564684684686u,0 2649.1330085085083u,0 2649.1340085085085u,1.5 2650.1105485485486u,1.5 2650.111548548549u,0 2652.065628628629u,0 2652.066628628629u,1.5 2653.0431686686684u,1.5 2653.0441686686686u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2673.5715095095093u,1.5 2673.5725095095095u,0 2674.5490495495496u,0 2674.55004954955u,1.5 2676.50412962963u,1.5 2676.50512962963u,0 2686.27953003003u,0 2686.28053003003u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2698.0100105105103u,1.5 2698.0110105105105u,0 2698.9875505505506u,0 2698.988550550551u,1.5 2699.9650905905905u,1.5 2699.9660905905907u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2708.7629509509507u,1.5 2708.763950950951u,0 2709.740490990991u,0 2709.741490990991u,1.5 2716.583271271271u,1.5 2716.584271271271u,0 2718.538351351351u,0 2718.5393513513513u,1.5 2719.5158913913915u,1.5 2719.5168913913917u,0 2721.4709714714713u,0 2721.4719714714715u,1.5 2722.4485115115112u,1.5 2722.4495115115114u,0 2726.3586716716713u,0 2726.3596716716715u,1.5 2727.3362117117117u,1.5 2727.337211711712u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2731.2463718718714u,0 2731.2473718718716u,1.5 2735.156532032032u,1.5 2735.157532032032u,0 2736.134072072072u,0 2736.135072072072u,1.5 2739.066692192192u,1.5 2739.067692192192u,0 2740.0442322322324u,0 2740.0452322322326u,1.5 2741.021772272272u,1.5 2741.022772272272u,0 2749.819632632633u,0 2749.820632632633u,1.5 2758.617492992993u,1.5 2758.618492992993u,0 2759.595033033033u,0 2759.596033033033u,1.5 2760.572573073073u,1.5 2760.573573073073u,0 2763.505193193193u,0 2763.506193193193u,1.5 2764.4827332332334u,1.5 2764.4837332332336u,0 2768.3928933933935u,0 2768.3938933933937u,1.5 2769.3704334334334u,1.5 2769.3714334334336u,0 2770.3479734734733u,0 2770.3489734734735u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2782.0784539539536u,1.5 2782.079453953954u,0 2790.876314314314u,0 2790.8773143143144u,1.5 2791.853854354354u,1.5 2791.8548543543543u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2793.8089344344344u,1.5 2793.8099344344346u,0 2794.7864744744743u,0 2794.7874744744745u,1.5 2804.561874874875u,1.5 2804.562874874875u,0 2814.337275275275u,0 2814.338275275275u,1.5 2821.1800555555556u,1.5 2821.1810555555558u,0 2822.1575955955955u,0 2822.1585955955957u,1.5 2828.022835835836u,1.5 2828.023835835836u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2846.5960965965965u,1.5 2846.5970965965967u,0 2847.573636636637u,0 2847.574636636637u,1.5 2848.5511766766763u,1.5 2848.5521766766765u,0 2849.5287167167166u,0 2849.529716716717u,1.5 2850.5062567567566u,1.5 2850.5072567567568u,0 2851.483796796797u,0 2851.484796796797u,1.5 2852.461336836837u,1.5 2852.462336836837u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2864.191817317317u,0 2864.1928173173173u,1.5 2876.899837837838u,1.5 2876.900837837838u,0 2877.877377877878u,0 2877.8783778778784u,1.5 2878.8549179179176u,1.5 2878.855917917918u,0 2880.809997997998u,0 2880.810997997998u,1.5 2881.787538038038u,1.5 2881.788538038038u,0 2882.765078078078u,0 2882.7660780780784u,1.5 2883.7426181181177u,1.5 2883.743618118118u,0 2889.607858358358u,0 2889.6088583583582u,1.5 2890.5853983983984u,1.5 2890.5863983983986u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2897.4281786786787u,1.5 2897.429178678679u,0 2898.4057187187186u,0 2898.406718718719u,1.5 2907.203579079079u,1.5 2907.2045790790794u,0 2908.1811191191186u,0 2908.182119119119u,1.5 2911.1137392392393u,1.5 2911.1147392392395u,0 2912.091279279279u,0 2912.0922792792794u,1.5 2913.068819319319u,1.5 2913.0698193193193u,0 2918.9340595595595u,0 2918.9350595595597u,1.5 2919.9115995995994u,1.5 2919.9125995995996u,0 2928.70945995996u,0 2928.71045995996u,1.5 2929.687u,1.5 2929.688u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2936.52978028028u,1.5 2936.5307802802804u,0 2937.50732032032u,0 2937.5083203203203u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2942.39502052052u,1.5 2942.3960205205203u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 2956.080581081081u,1.5 2956.0815810810814u,0 2957.0581211211206u,0 2957.059121121121u,1.5 2960.968281281281u,1.5 2960.9692812812814u,0 2961.945821321321u,0 2961.9468213213213u,1.5 2962.923361361361u,1.5 2962.924361361361u,0 2964.8784414414413u,0 2964.8794414414415u,1.5 2965.8559814814816u,1.5 2965.856981481482u,0 2966.833521521521u,0 2966.8345215215213u,1.5 2967.8110615615615u,1.5 2967.8120615615617u,0 2968.7886016016014u,0 2968.7896016016016u,1.5 2969.7661416416418u,1.5 2969.767141641642u,0 2970.7436816816817u,0 2970.744681681682u,1.5 2972.6987617617615u,1.5 2972.6997617617617u,0 2974.6538418418418u,0 2974.654841841842u,1.5 2975.631381881882u,1.5 2975.6323818818823u,0 2980.519082082082u,0 2980.5200820820824u,1.5 2981.4966221221216u,1.5 2981.497622122122u,0 2983.451702202202u,0 2983.452702202202u,1.5 2984.4292422422423u,1.5 2984.4302422422425u,0 2986.384322322322u,0 2986.3853223223223u,1.5 2987.361862362362u,1.5 2987.362862362362u,0 2989.3169424424423u,0 2989.3179424424425u,1.5 2990.2944824824826u,1.5 2990.295482482483u,0 2993.2271026026024u,0 2993.2281026026026u,1.5 2994.2046426426427u,1.5 2994.205642642643u,0 2999.0923428428428u,0 2999.093342842843u,1.5 3000.069882882883u,1.5 3000.0708828828833u,0 3003.980043043043u,0 3003.9810430430434u,1.5 3004.957583083083u,1.5 3004.9585830830833u,0 3010.822823323323u,0 3010.8238233233233u,1.5 3011.800363363363u,1.5 3011.801363363363u,0 3014.7329834834836u,0 3014.733983483484u,1.5 3015.710523523523u,1.5 3015.7115235235233u,0 3017.6656036036034u,0 3017.6666036036036u,1.5 3018.6431436436437u,1.5 3018.644143643644u,0 3022.553303803804u,0 3022.554303803804u,1.5 3023.5308438438437u,1.5 3023.531843843844u,0 3026.463463963964u,0 3026.464463963964u,1.5 3027.441004004004u,1.5 3027.442004004004u,0 3028.418544044044u,0 3028.4195440440444u,1.5 3029.396084084084u,1.5 3029.3970840840843u,0 3030.373624124124u,0 3030.3746241241242u,1.5 3032.328704204204u,1.5 3032.329704204204u,0 3033.306244244244u,0 3033.3072442442444u,1.5 3036.238864364364u,1.5 3036.239864364364u,0 3037.2164044044043u,0 3037.2174044044045u,1.5 3039.1714844844846u,1.5 3039.172484484485u,0 3040.149024524524u,0 3040.1500245245243u,1.5 3060.677365365365u,1.5 3060.678365365365u,0 3061.6549054054053u,0 3061.6559054054055u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3064.587525525525u,0 3064.5885255255253u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3069.4752257257255u,0 3069.4762257257257u,1.5 3070.4527657657654u,1.5 3070.4537657657656u,0 3074.3629259259255u,0 3074.3639259259257u,1.5 3075.340465965966u,1.5 3075.341465965966u,0 3085.115866366366u,0 3085.116866366366u,1.5 3086.0934064064063u,1.5 3086.0944064064065u,0 3089.026026526526u,0 3089.0270265265262u,1.5 3098.8014269269265u,1.5 3098.8024269269267u,0 3099.778966966967u,0 3099.779966966967u,1.5 3102.711587087087u,1.5 3102.7125870870873u,0 3103.689127127127u,0 3103.690127127127u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3108.576827327327u,0 3108.577827327327u,1.5 3109.554367367367u,1.5 3109.555367367367u,0 3120.307307807808u,0 3120.308307807808u,1.5 3121.2848478478477u,1.5 3121.285847847848u,0 3122.262387887888u,0 3122.2633878878883u,1.5 3132.037788288288u,1.5 3132.0387882882883u,0 3133.0153283283285u,0 3133.0163283283287u,1.5 3134.9704084084083u,1.5 3134.9714084084085u,0 3136.9254884884886u,0 3136.9264884884888u,1.5 3137.9030285285285u,1.5 3137.9040285285287u,0 3145.7233488488487u,0 3145.724348848849u,1.5 3146.700888888889u,1.5 3146.7018888888892u,0 3147.678428928929u,0 3147.679428928929u,1.5 3148.655968968969u,1.5 3148.656968968969u,0 3149.633509009009u,0 3149.634509009009u,1.5 3151.588589089089u,1.5 3151.5895890890893u,0 3152.5661291291294u,0 3152.5671291291296u,1.5 3161.3639894894895u,1.5 3161.3649894894897u,0 3162.3415295295295u,0 3162.3425295295297u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3164.2966096096093u,0 3164.2976096096095u,1.5 3165.2741496496496u,1.5 3165.27514964965u,0 3174.0720100100098u,0 3174.07301001001u,1.5 3175.04955005005u,1.5 3175.0505500500503u,0 3176.02709009009u,0 3176.0280900900902u,1.5 3183.8474104104102u,1.5 3183.8484104104105u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3187.7575705705704u,1.5 3187.7585705705706u,0 3195.577890890891u,0 3195.578890890891u,1.5 3196.555430930931u,1.5 3196.556430930931u,0 3197.532970970971u,0 3197.533970970971u,1.5 3209.263451451451u,1.5 3209.2644514514514u,0 3216.106231731732u,0 3216.107231731732u,1.5 3217.0837717717714u,1.5 3217.0847717717716u,0 3218.0613118118117u,0 3218.062311811812u,1.5 3219.0388518518516u,1.5 3219.039851851852u,0 3220.016391891892u,0 3220.017391891892u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3238.5896526526526u,0 3238.590652652653u,1.5 3240.544732732733u,1.5 3240.545732732733u,0 3241.5222727727723u,0 3241.5232727727725u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3261.0730735735733u,0 3261.0740735735735u,1.5 3262.050613613613u,1.5 3262.0516136136134u,0 3263.0281536536536u,0 3263.029153653654u,1.5 3269.870933933934u,1.5 3269.871933933934u,0 3270.848473973974u,0 3270.849473973974u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3273.781094094094u,1.5 3273.782094094094u,0 3280.6238743743743u,0 3280.6248743743745u,1.5 3281.601414414414u,1.5 3281.6024144144144u,0 3283.5564944944945u,0 3283.5574944944947u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3301.152215215215u,0 3301.1532152152154u,1.5 3302.129755255255u,1.5 3302.1307552552553u,0 3303.1072952952954u,0 3303.1082952952956u,1.5 3306.039915415415u,1.5 3306.0409154154154u,0 3307.017455455455u,0 3307.0184554554553u,1.5 3312.8826956956955u,1.5 3312.8836956956957u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3315.8153158158157u,1.5 3315.816315815816u,0 3317.770395895896u,0 3317.771395895896u,1.5 3318.747935935936u,1.5 3318.748935935936u,0 3325.590716216216u,0 3325.5917162162164u,1.5 3326.568256256256u,1.5 3326.5692562562563u,0 3327.5457962962964u,0 3327.5467962962966u,1.5 3328.5233363363363u,1.5 3328.5243363363365u,0 3329.5008763763763u,0 3329.5018763763765u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3337.3211966966965u,0 3337.3221966966967u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3350.029217217217u,0 3350.0302172172173u,1.5 3351.006757257257u,1.5 3351.0077572572573u,0 3351.9842972972974u,0 3351.9852972972976u,1.5 3361.7596976976974u,1.5 3361.7606976976977u,0 3363.7147777777773u,0 3363.7157777777775u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3379.355418418418u,0 3379.3564184184183u,1.5 3382.2880385385383u,1.5 3382.2890385385385u,0 3383.2655785785787u,0 3383.266578578579u,1.5 3388.1532787787787u,1.5 3388.154278778779u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.0185190190186u,0 3394.019519019019u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3398.906219219219u,0 3398.9072192192193u,1.5 3399.883759259259u,1.5 3399.884759259259u,0 3408.681619619619u,0 3408.6826196196193u,1.5 3409.6591596596595u,1.5 3409.6601596596597u,0 3410.6366996996994u,0 3410.6376996996996u,1.5 3411.61423973974u,1.5 3411.61523973974u,0 3412.5917797797797u,0 3412.59277977978u,1.5 3414.5468598598595u,1.5 3414.5478598598597u,0 3415.5243998999u,0 3415.5253998999u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3437.0302807807807u,1.5 3437.031280780781u,0 3438.0078208208206u,0 3438.008820820821u,1.5 3438.9853608608605u,1.5 3438.9863608608607u,0 3460.4912417417418u,0 3460.492241741742u,1.5 3461.4687817817817u,1.5 3461.469781781782u,0 3465.378941941942u,0 3465.379941941942u,1.5 3466.356481981982u,1.5 3466.3574819819823u,0 3467.3340220220216u,0 3467.335022022022u,1.5 3468.311562062062u,1.5 3468.312562062062u,0 3469.289102102102u,0 3469.290102102102u,1.5 3470.2666421421422u,1.5 3470.2676421421424u,0 3472.221722222222u,0 3472.2227222222223u,1.5 3473.199262262262u,1.5 3473.200262262262u,0 3474.1768023023023u,0 3474.1778023023026u,1.5 3475.1543423423423u,1.5 3475.1553423423425u,0 3476.1318823823826u,0 3476.132882382383u,1.5 3478.0869624624625u,1.5 3478.0879624624627u,0 3479.0645025025024u,0 3479.0655025025026u,1.5 3481.0195825825826u,1.5 3481.020582582583u,0 3481.997122622622u,0 3481.9981226226223u,1.5 3482.9746626626625u,1.5 3482.9756626626627u,0 3483.9522027027024u,0 3483.9532027027026u,1.5 3493.727603103103u,1.5 3493.728603103103u,0 3494.7051431431432u,0 3494.7061431431434u,1.5 3501.547923423423u,1.5 3501.5489234234233u,0 3502.5254634634634u,0 3502.5264634634636u,1.5 3521.098724224224u,1.5 3521.0997242242242u,0 3522.076264264264u,0 3522.077264264264u,1.5 3525.0088843843846u,1.5 3525.009884384385u,0 3526.9639644644644u,0 3526.9649644644646u,1.5 3527.9415045045043u,1.5 3527.9425045045045u,0 3529.8965845845846u,0 3529.897584584585u,1.5 3530.8741246246245u,1.5 3530.8751246246247u,0 3531.8516646646644u,0 3531.8526646646646u,1.5 3533.8067447447447u,1.5 3533.807744744745u,0 3535.7618248248245u,0 3535.7628248248247u,1.5 3536.7393648648645u,1.5 3536.7403648648647u,0 3537.716904904905u,0 3537.717904904905u,1.5 3538.6944449449447u,1.5 3538.695444944945u,0 3540.6495250250246u,0 3540.6505250250248u,1.5 3541.627065065065u,1.5 3541.628065065065u,0 3561.1778658658654u,0 3561.1788658658656u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3564.110485985986u,0 3564.1114859859863u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.998186186186u,1.5 3568.9991861861863u,0 3569.975726226226u,0 3569.976726226226u,1.5 3583.6612867867866u,1.5 3583.662286786787u,0 3584.6388268268265u,0 3584.6398268268267u,1.5 3586.593906906907u,1.5 3586.594906906907u,0 3588.548986986987u,0 3588.5499869869873u,1.5 3589.5265270270265u,1.5 3589.5275270270267u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3609.0773278278275u,0 3609.0783278278277u,1.5 3618.852728228228u,1.5 3618.853728228228u,0 3619.830268268268u,0 3619.831268268268u,1.5 3621.785348348348u,1.5 3621.7863483483484u,0 3622.7628883883885u,0 3622.7638883883888u,1.5 3623.740428428428u,1.5 3623.741428428428u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3650.1340095095093u,1.5 3650.1350095095095u,0 3651.1115495495496u,0 3651.11254954955u,1.5 3652.0890895895895u,1.5 3652.0900895895898u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3669.6848103103102u,1.5 3669.6858103103104u,0 3670.66235035035u,0 3670.6633503503504u,1.5 3675.5500505505506u,1.5 3675.551050550551u,0 3676.5275905905905u,0 3676.5285905905907u,1.5 3677.505130630631u,1.5 3677.506130630631u,0 3681.4152907907906u,0 3681.4162907907908u,1.5 3682.392830830831u,1.5 3682.393830830831u,0 3685.3254509509507u,0 3685.326450950951u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3697.0559314314314u,1.5 3697.0569314314316u,0 3698.0334714714713u,0 3698.0344714714715u,1.5 3699.0110115115112u,1.5 3699.0120115115114u,0 3704.8762517517516u,0 3704.877251751752u,1.5 3705.8537917917915u,1.5 3705.8547917917917u,0 3707.8088718718714u,0 3707.8098718718716u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3718.561812312312u,1.5 3718.5628123123124u,0 3719.539352352352u,0 3719.5403523523523u,1.5 3720.5168923923925u,1.5 3720.5178923923927u,0 3728.3372127127127u,0 3728.338212712713u,1.5 3729.3147527527526u,1.5 3729.315752752753u,0 3730.292292792793u,0 3730.293292792793u,1.5 3733.2249129129127u,1.5 3733.225912912913u,0 3734.2024529529526u,0 3734.203452952953u,1.5 3740.067693193193u,1.5 3740.068693193193u,0 3746.9104734734733u,0 3746.9114734734735u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3758.6409539539536u,1.5 3758.641953953954u,0 3759.618493993994u,0 3759.619493993994u,1.5 3760.596034034034u,1.5 3760.597034034034u,0 3762.5511141141137u,0 3762.552114114114u,1.5 3763.528654154154u,1.5 3763.5296541541543u,0 3770.3714344344344u,0 3770.3724344344346u,1.5 3780.146834834835u,1.5 3780.147834834835u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3800.6751756756753u,1.5 3800.6761756756755u,0 3801.6527157157157u,0 3801.653715715716u,1.5 3804.585335835836u,1.5 3804.586335835836u,0 3815.338276276276u,0 3815.339276276276u,1.5 3829.023836836837u,1.5 3829.024836836837u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3851.5072577577575u,1.5 3851.5082577577577u,0 3862.260198198198u,0 3862.261198198198u,1.5 3864.2152782782778u,1.5 3864.216278278278u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3873.013138638639u,1.5 3873.014138638639u,0 3873.9906786786783u,0 3873.9916786786785u,1.5 3877.900838838839u,1.5 3877.901838838839u,0 3878.878378878879u,0 3878.8793788788794u,1.5 3879.8559189189186u,1.5 3879.856918918919u,0 3889.631319319319u,0 3889.6323193193193u,1.5 3890.608859359359u,1.5 3890.6098593593592u,0 3892.5639394394393u,0 3892.5649394394395u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3907.22704004004u,1.5 3907.22804004004u,0 3908.20458008008u,0 3908.2055800800804u,1.5 3909.1821201201196u,1.5 3909.18312012012u,0 3910.1596601601605u,0 3910.1606601601607u,1.5 3913.09228028028u,1.5 3913.0932802802804u,0 3929.710460960961u,0 3929.711460960961u,1.5 3930.688001001001u,1.5 3930.689001001001u,0 3931.665541041041u,0 3931.666541041041u,1.5 3932.643081081081u,1.5 3932.6440810810814u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3937.530781281281u,0 3937.5317812812814u,1.5 3958.0591221221216u,1.5 3958.060122122122u,0 3959.0366621621624u,0 3959.0376621621626u,1.5 3964.9019024024024u,1.5 3964.9029024024026u,0 3965.879442442442u,0 3965.880442442442u,1.5 3967.834522522522u,1.5 3967.8355225225223u,0 3969.7896026026024u,0 3969.7906026026026u,1.5 3970.7671426426423u,1.5 3970.7681426426425u,0 3971.7446826826827u,0 3971.745682682683u,1.5 3972.7222227227226u,1.5 3972.7232227227228u,0 3974.677302802803u,0 3974.678302802803u,1.5 3976.632382882883u,1.5 3976.6333828828833u,0 3977.6099229229226u,0 3977.610922922923u,1.5 3978.5874629629634u,1.5 3978.5884629629636u,0 3985.430243243243u,0 3985.431243243243u,1.5 3986.407783283283u,1.5 3986.4087832832834u,0 3990.317943443443u,0 3990.318943443443u,1.5 3991.2954834834836u,1.5 3991.296483483484u,0 3994.2281036036034u,0 3994.2291036036036u,1.5 3995.2056436436433u,1.5 3995.2066436436435u,0 3998.138263763764u,0 3998.139263763764u,1.5 3999.115803803804u,1.5 3999.116803803804u,0 4004.9810440440438u,0 4004.982044044044u,1.5 4005.958584084084u,1.5 4005.9595840840843u,0 4010.846284284284u,0 4010.8472842842843u,1.5 4011.823824324324u,1.5 4011.8248243243243u,0 4012.8013643643644u,0 4012.8023643643646u,1.5 4013.7789044044043u,1.5 4013.7799044044045u,0 4018.6666046046043u,0 4018.6676046046045u,1.5 4019.6441446446443u,1.5 4019.6451446446445u,0 4023.554304804805u,0 4023.555304804805u,1.5 4024.5318448448443u,1.5 4024.5328448448445u,0 4025.509384884885u,0 4025.5103848848853u,1.5 4026.4869249249246u,1.5 4026.4879249249248u,0 4027.4644649649654u,0 4027.4654649649656u,1.5 4028.442005005005u,1.5 4028.443005005005u,0 4029.4195450450447u,0 4029.420545045045u,1.5 4031.374625125125u,1.5 4031.375625125125u,0 4032.3521651651654u,0 4032.3531651651656u,1.5 4033.329705205205u,1.5 4033.330705205205u,0 4035.284785285285u,0 4035.2857852852853u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4069.4986866866866u,1.5 4069.499686686687u,0 4070.4762267267265u,0 4070.4772267267267u,1.5 4071.453766766767u,1.5 4071.454766766767u,0 4078.2965470470467u,0 4078.297547047047u,1.5 4079.274087087087u,1.5 4079.2750870870873u,0 4081.2291671671674u,0 4081.2301671671676u,1.5 4082.206707207207u,1.5 4082.207707207207u,0 4087.0944074074073u,0 4087.0954074074075u,1.5 4089.0494874874876u,1.5 4089.0504874874878u,0 4090.027027527527u,0 4090.0280275275272u,1.5 4093.9371876876876u,1.5 4093.938187687688u,0 4094.9147277277275u,0 4094.9157277277277u,1.5 4103.7125880880885u,1.5 4103.713588088089u,0 4104.690128128128u,0 4104.691128128128u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4120.330768768769u,0 4120.3317687687695u,1.5 4121.308308808809u,1.5 4121.309308808809u,0 4122.285848848848u,0 4122.286848848848u,1.5 4124.240928928929u,1.5 4124.241928928929u,0 4125.218468968969u,0 4125.2194689689695u,1.5 4131.083709209209u,1.5 4131.084709209209u,0 4132.061249249249u,0 4132.062249249249u,1.5 4136.948949449449u,1.5 4136.949949449449u,0 4138.904029529529u,0 4138.905029529529u,1.5 4139.881569569569u,1.5 4139.88256956957u,0 4148.67942992993u,0 4148.68042992993u,1.5 4149.65696996997u,1.5 4149.6579699699705u,0 4150.63451001001u,0 4150.63551001001u,1.5 4160.40991041041u,1.5 4160.41091041041u,0 4161.38745045045u,0 4161.38845045045u,1.5 4162.3649904904905u,1.5 4162.365990490491u,0 4164.32007057057u,0 4164.321070570571u,1.5 4165.297610610611u,1.5 4165.298610610611u,0 4172.140390890891u,0 4172.141390890891u,1.5 4173.117930930931u,1.5 4173.118930930931u,0 4174.095470970971u,0 4174.0964709709715u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4187.781031531531u,1.5 4187.782031531531u,0 4193.646271771772u,0 4193.6472717717725u,1.5 4194.623811811812u,1.5 4194.624811811812u,0 4197.556431931932u,0 4197.557431931932u,1.5 4198.533971971972u,1.5 4198.5349719719725u,0 4199.511512012012u,0 4199.512512012012u,1.5 4206.3542922922925u,1.5 4206.355292292293u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4210.264452452452u,0 4210.265452452452u,1.5 4211.2419924924925u,1.5 4211.242992492493u,0 4217.107232732732u,0 4217.108232732732u,1.5 4218.084772772773u,1.5 4218.085772772773u,0 4219.062312812813u,0 4219.063312812813u,1.5 4228.837713213213u,1.5 4228.838713213213u,0 4230.7927932932935u,0 4230.793793293294u,1.5 4231.770333333333u,1.5 4231.771333333333u,0 4237.635573573573u,0 4237.6365735735735u,1.5 4238.613113613614u,1.5 4238.614113613614u,0 4240.5681936936935u,0 4240.569193693694u,1.5 4243.500813813814u,1.5 4243.501813813814u,0 4244.478353853853u,0 4244.479353853853u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4261.096534534534u,0 4261.097534534534u,1.5 4263.051614614615u,1.5 4263.052614614615u,0 4264.029154654655u,0 4264.030154654655u,1.5 4266.961774774775u,1.5 4266.962774774775u,0 4267.939314814815u,0 4267.940314814815u,1.5 4271.849474974975u,1.5 4271.850474974975u,0 4279.669795295295u,0 4279.670795295296u,1.5 4280.647335335335u,1.5 4280.648335335335u,0 4281.624875375375u,0 4281.6258753753755u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4301.175676176176u,0 4301.176676176176u,1.5 4302.153216216216u,1.5 4302.154216216216u,0 4303.130756256257u,0 4303.131756256257u,1.5 4315.838776776777u,1.5 4315.839776776777u,0 4316.816316816817u,0 4316.817316816817u,1.5 4317.793856856857u,1.5 4317.794856856857u,0 4325.614177177177u,0 4325.615177177177u,1.5 4326.591717217217u,1.5 4326.592717217217u,0 4327.569257257258u,0 4327.570257257258u,1.5 4328.546797297297u,1.5 4328.547797297298u,0 4329.524337337337u,0 4329.525337337337u,1.5 4334.412037537537u,1.5 4334.413037537537u,0 4335.389577577577u,0 4335.3905775775775u,1.5 4338.322197697697u,1.5 4338.323197697698u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4351.030218218218u,0 4351.031218218218u,1.5 4352.007758258259u,1.5 4352.008758258259u,0 4352.985298298298u,0 4352.986298298299u,1.5 4360.805618618619u,1.5 4360.806618618619u,0 4361.783158658659u,0 4361.784158658659u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4376.44625925926u,0 4376.44725925926u,1.5 4377.423799299299u,1.5 4377.4247992993u,0 4379.378879379379u,0 4379.379879379379u,1.5 4392.086899899899u,1.5 4392.0878998999u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.01952002002u,0 4395.02052002002u,1.5 4396.9746001001u,1.5 4396.975600100101u,0 4407.72754054054u,0 4407.72854054054u,1.5 4408.70508058058u,1.5 4408.70608058058u,0 4409.682620620621u,0 4409.683620620621u,1.5 4410.660160660661u,1.5 4410.661160660661u,0 4412.61524074074u,0 4412.61624074074u,1.5 4414.570320820821u,1.5 4414.571320820821u,0 4415.547860860861u,0 4415.548860860861u,1.5 4430.210961461462u,1.5 4430.211961461462u,0 4431.188501501501u,0 4431.189501501502u,1.5 4432.166041541541u,1.5 4432.167041541541u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4439.008821821822u,0 4439.009821821822u,1.5 4439.986361861862u,1.5 4439.987361861862u,0 4440.963901901901u,0 4440.964901901902u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4457.582082582582u,0 4457.583082582582u,1.5 4458.559622622623u,1.5 4458.560622622623u,0 4459.537162662663u,0 4459.538162662663u,1.5 4460.514702702702u,1.5 4460.515702702703u,0 4467.357482982983u,0 4467.358482982983u,1.5 4468.335023023023u,1.5 4468.336023023023u,0 4469.312563063063u,0 4469.313563063063u,1.5 4471.267643143143u,1.5 4471.268643143143u,0 4472.245183183183u,0 4472.246183183183u,1.5 4473.222723223223u,1.5 4473.223723223223u,0 4474.200263263264u,0 4474.201263263264u,1.5 4475.177803303303u,1.5 4475.1788033033035u,0 4476.155343343343u,0 4476.156343343343u,1.5 4478.1104234234235u,1.5 4478.111423423424u,0 4479.087963463464u,0 4479.088963463464u,1.5 4482.9981236236235u,1.5 4482.999123623624u,0 4483.975663663664u,0 4483.976663663664u,1.5 4484.953203703703u,1.5 4484.954203703704u,0 4485.930743743743u,0 4485.931743743743u,1.5 4491.795983983984u,1.5 4491.796983983984u,0 4492.773524024024u,0 4492.774524024024u,1.5 4494.728604104104u,1.5 4494.7296041041045u,0 4495.706144144144u,0 4495.707144144144u,1.5 4503.526464464465u,1.5 4503.527464464465u,0 4504.504004504504u,0 4504.5050045045045u,1.5 4506.459084584585u,1.5 4506.460084584585u,0 4507.4366246246245u,0 4507.437624624625u,1.5 4510.369244744744u,1.5 4510.370244744744u,0 4511.346784784785u,0 4511.347784784785u,1.5 4514.279404904904u,1.5 4514.280404904905u,0 4515.256944944945u,0 4515.257944944945u,1.5 4519.167105105105u,1.5 4519.1681051051055u,0 4520.144645145145u,0 4520.145645145145u,1.5 4522.099725225225u,1.5 4522.100725225225u,0 4523.077265265266u,0 4523.078265265266u,1.5 4525.032345345345u,1.5 4525.033345345345u,0 4526.9874254254255u,0 4526.988425425426u,1.5 4528.942505505505u,1.5 4528.9435055055055u,0 4529.920045545545u,0 4529.921045545545u,1.5 4531.8751256256255u,1.5 4531.876125625626u,0 4536.7628258258255u,0 4536.763825825826u,1.5 4537.740365865866u,1.5 4537.741365865866u,0 4539.695445945946u,0 4539.696445945946u,1.5 4540.672985985986u,1.5 4540.673985985986u,0 4542.628066066066u,0 4542.629066066066u,1.5 4543.605606106106u,1.5 4543.6066061061065u,0 4562.178866866867u,0 4562.179866866867u,1.5 4563.156406906906u,1.5 4563.1574069069065u,0 4565.111486986987u,0 4565.112486986987u,1.5 4569.021647147147u,1.5 4569.022647147147u,0 4569.999187187187u,0 4570.000187187187u,1.5 4584.662287787788u,1.5 4584.663287787788u,0 4585.6398278278275u,0 4585.640827827828u,1.5 4586.617367867868u,1.5 4586.618367867868u,0 4587.594907907907u,0 4587.5959079079075u,1.5 4588.572447947948u,1.5 4588.573447947948u,0 4590.5275280280275u,0 4590.528528028028u,1.5 4591.505068068068u,1.5 4591.506068068068u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4607.145708708708u,1.5 4607.1467087087085u,0 4608.123248748749u,0 4608.124248748749u,1.5 4620.83126926927u,1.5 4620.83226926927u,0 4622.786349349349u,0 4622.787349349349u,1.5 4623.763889389389u,1.5 4623.764889389389u,0 4634.5168298298295u,0 4634.51782982983u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4637.44944994995u,0 4637.45044994995u,1.5 4640.38207007007u,1.5 4640.38307007007u,0 4641.35961011011u,0 4641.36061011011u,1.5 4649.17993043043u,1.5 4649.180930430431u,0 4651.13501051051u,0 4651.1360105105105u,1.5 4652.11255055055u,1.5 4652.11355055055u,0 4653.090090590591u,0 4653.091090590591u,1.5 4654.06763063063u,1.5 4654.068630630631u,0 4659.932870870871u,0 4659.933870870871u,1.5 4660.91041091091u,1.5 4660.9114109109105u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4666.775651151151u,1.5 4666.776651151151u,0 4667.753191191191u,0 4667.754191191191u,1.5 4671.663351351351u,1.5 4671.664351351351u,0 4672.640891391391u,0 4672.641891391391u,1.5 4673.618431431431u,1.5 4673.619431431432u,0 4685.348911911911u,0 4685.3499119119115u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4687.303991991992u,0 4687.304991991992u,1.5 4688.2815320320315u,1.5 4688.282532032032u,0 4689.259072072072u,0 4689.260072072072u,1.5 4697.079392392392u,1.5 4697.080392392392u,0 4698.056932432432u,0 4698.057932432433u,1.5 4699.034472472473u,1.5 4699.035472472473u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4709.787412912912u,0 4709.7884129129125u,1.5 4718.585273273274u,1.5 4718.586273273274u,0 4720.540353353353u,0 4720.541353353353u,1.5 4721.517893393393u,1.5 4721.518893393393u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4740.091154154154u,1.5 4740.092154154154u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 4760.619494994995u,1.5 4760.620494994995u,0 4761.597035035034u,0 4761.598035035035u,1.5 4762.574575075075u,1.5 4762.575575075075u,0 4770.394895395395u,0 4770.395895395395u,1.5 4772.349975475476u,1.5 4772.350975475476u,0 4773.327515515515u,0 4773.328515515515u,1.5 4777.237675675676u,1.5 4777.238675675676u,0 4778.215215715715u,0 4778.216215715715u,1.5 4781.147835835835u,1.5 4781.148835835836u,0 4784.0804559559565u,0 4784.081455955957u,1.5 4785.057995995996u,1.5 4785.058995995996u,0 4792.878316316316u,0 4792.879316316316u,1.5 4795.810936436436u,1.5 4795.811936436437u,0 4796.788476476477u,0 4796.789476476477u,1.5 4804.608796796797u,1.5 4804.609796796797u,0 4815.361737237236u,0 4815.362737237237u,1.5 4816.339277277278u,1.5 4816.340277277278u,0 4817.316817317317u,0 4817.317817317317u,1.5 4823.1820575575575u,1.5 4823.183057557558u,0 4824.159597597598u,0 4824.160597597598u,1.5 4825.137137637637u,1.5 4825.138137637638u,0 4826.114677677678u,0 4826.115677677678u,1.5 4827.092217717717u,1.5 4827.093217717717u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4849.575638638638u,1.5 4849.5766386386385u,0 4850.553178678679u,0 4850.554178678679u,1.5 4851.530718718718u,1.5 4851.531718718718u,0 4852.508258758759u,0 4852.50925875876u,1.5 4853.485798798799u,1.5 4853.486798798799u,0 4865.21627927928u,0 4865.21727927928u,1.5 4876.94675975976u,1.5 4876.947759759761u,0 4877.9242997998u,0 4877.9252997998u,1.5 4878.901839839839u,1.5 4878.9028398398395u,0 4879.87937987988u,0 4879.88037987988u,1.5 4880.85691991992u,1.5 4880.85791991992u,0 4882.812u,0 4882.813u,1.5 4883.789540040039u,1.5 4883.79054004004u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4895.52002052052u,1.5 4895.52102052052u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4907.250501001001u,1.5 4907.251501001001u,0 4908.22804104104u,0 4908.229041041041u,1.5 4911.160661161161u,1.5 4911.161661161162u,0 4912.138201201201u,0 4912.139201201201u,1.5 4914.093281281282u,1.5 4914.094281281282u,0 4917.025901401401u,0 4917.026901401401u,1.5 4918.003441441441u,1.5 4918.0044414414415u,0 4930.711461961962u,0 4930.712461961963u,1.5 4931.689002002002u,1.5 4931.690002002002u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4935.599162162162u,0 4935.600162162163u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4939.509322322322u,1.5 4939.510322322322u,0 4940.486862362362u,0 4940.487862362363u,1.5 4964.925363363363u,1.5 4964.926363363364u,0 4965.902903403403u,0 4965.903903403403u,1.5 4969.813063563563u,1.5 4969.814063563564u,0 4970.790603603604u,0 4970.791603603604u,1.5 4971.768143643643u,1.5 4971.7691436436435u,0 4972.745683683684u,0 4972.746683683684u,1.5 4973.723223723723u,1.5 4973.724223723723u,0 4974.700763763764u,0 4974.701763763765u,1.5 4976.655843843843u,1.5 4976.6568438438435u,0 4977.633383883884u,0 4977.634383883884u,1.5 4978.610923923924u,1.5 4978.611923923924u,0 4983.498624124124u,0 4983.499624124124u,1.5 4984.476164164164u,1.5 4984.477164164165u,0 4988.386324324324u,0 4988.387324324324u,1.5 4989.363864364364u,1.5 4989.364864364365u,0 5003.049424924925u,0 5003.050424924925u,1.5 5004.026964964965u,1.5 5004.027964964966u,0 5005.982045045044u,0 5005.9830450450445u,1.5 5006.959585085086u,1.5 5006.960585085086u,0 5014.779905405405u,0 5014.780905405405u,1.5 5015.757445445445u,1.5 5015.758445445445u,0 5017.712525525525u,0 5017.713525525525u,1.5 5018.690065565565u,1.5 5018.691065565566u,0 5020.645145645645u,0 5020.646145645645u,1.5 5021.622685685686u,1.5 5021.623685685686u,0 5022.600225725725u,0 5022.601225725725u,1.5 5024.555305805806u,1.5 5024.556305805806u,0 5025.532845845845u,0 5025.5338458458455u,1.5 5026.510385885886u,1.5 5026.511385885886u,0 5028.465465965966u,0 5028.466465965967u,1.5 5029.443006006006u,1.5 5029.444006006006u,0 5031.398086086087u,0 5031.399086086087u,1.5 5033.353166166166u,1.5 5033.354166166167u,0 5034.330706206206u,0 5034.331706206206u,1.5 5042.151026526526u,1.5 5042.152026526526u,0 5043.128566566566u,0 5043.129566566567u,1.5 5055.8365870870875u,1.5 5055.837587087088u,0 5056.814127127127u,0 5056.815127127127u,1.5 5059.746747247247u,1.5 5059.747747247247u,0 5060.724287287288u,0 5060.725287287288u,1.5 5061.701827327327u,1.5 5061.702827327327u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5067.567067567567u,0 5067.568067567568u,1.5 5068.544607607608u,1.5 5068.545607607608u,0 5071.477227727727u,0 5071.478227727727u,1.5 5072.454767767768u,1.5 5072.4557677677685u,0 5084.185248248248u,0 5084.186248248248u,1.5 5085.1627882882885u,1.5 5085.163788288289u,0 5087.117868368368u,0 5087.118868368369u,1.5 5088.095408408408u,1.5 5088.096408408408u,0 5089.072948448448u,0 5089.073948448448u,1.5 5092.983108608609u,1.5 5092.984108608609u,0 5093.960648648648u,0 5093.961648648648u,1.5 5095.915728728728u,1.5 5095.916728728728u,0 5096.893268768769u,0 5096.8942687687695u,1.5 5103.736049049048u,1.5 5103.737049049048u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5108.623749249249u,1.5 5108.624749249249u,0 5117.42160960961u,0 5117.42260960961u,1.5 5118.399149649649u,1.5 5118.400149649649u,0 5121.33176976977u,0 5121.3327697697705u,1.5 5122.30930980981u,1.5 5122.31030980981u,0 5123.286849849849u,0 5123.287849849849u,1.5 5134.0397902902905u,1.5 5134.040790290291u,0 5135.01733033033u,0 5135.01833033033u,1.5 5136.97241041041u,1.5 5136.97341041041u,0 5137.94995045045u,0 5137.95095045045u,1.5 5138.9274904904905u,1.5 5138.928490490491u,0 5148.702890890891u,0 5148.703890890891u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5163.3659914914915u,0 5163.366991491492u,1.5 5164.343531531531u,1.5 5164.344531531531u,0 5173.1413918918915u,0 5173.142391891892u,1.5 5174.118931931932u,1.5 5174.119931931932u,0 5175.096471971972u,0 5175.0974719719725u,1.5 5181.939252252252u,1.5 5181.940252252252u,0 5182.9167922922925u,0 5182.917792292293u,1.5 5185.849412412412u,1.5 5185.850412412412u,0 5186.826952452452u,0 5186.827952452452u,1.5 5187.8044924924925u,1.5 5187.805492492493u,0 5197.5798928928925u,0 5197.580892892893u,1.5 5207.3552932932935u,1.5 5207.356293293294u,0 5208.332833333333u,0 5208.333833333333u,1.5 5209.310373373373u,1.5 5209.3113733733735u,0 5210.287913413413u,0 5210.288913413413u,1.5 5211.265453453453u,1.5 5211.266453453453u,0 5217.1306936936935u,0 5217.131693693694u,1.5 5218.108233733733u,1.5 5218.109233733733u,0 5219.085773773774u,0 5219.086773773774u,1.5 5220.063313813814u,1.5 5220.064313813814u,0 5221.040853853853u,0 5221.041853853853u,1.5 5228.861174174174u,1.5 5228.8621741741745u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5239.614114614615u,0 5239.615114614615u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5257.209835335335u,0 5257.210835335335u,1.5 5258.187375375375u,1.5 5258.1883753753755u,0 5260.142455455456u,0 5260.143455455456u,1.5 5261.1199954954955u,1.5 5261.120995495496u,0 5262.097535535535u,0 5262.098535535535u,1.5 5264.052615615616u,1.5 5264.053615615616u,0 5265.030155655656u,0 5265.031155655656u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5274.805556056056u,0 5274.806556056056u,1.5 5275.783096096096u,1.5 5275.784096096097u,0 5281.648336336336u,0 5281.649336336336u,1.5 5282.625876376376u,1.5 5282.6268763763765u,0 5283.603416416417u,0 5283.604416416417u,1.5 5287.513576576576u,1.5 5287.5145765765765u,0 5288.491116616617u,0 5288.492116616617u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5303.154217217217u,0 5303.155217217217u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5316.839777777778u,1.5 5316.840777777778u,0 5327.592718218218u,0 5327.593718218218u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5346.165978978979u,0 5346.166978978979u,1.5 5347.143519019019u,1.5 5347.144519019019u,0 5349.098599099099u,0 5349.0995990991u,1.5 5350.076139139139u,1.5 5350.077139139139u,0 5352.031219219219u,0 5352.032219219219u,1.5 5359.851539539539u,1.5 5359.852539539539u,0 5360.829079579579u,0 5360.830079579579u,1.5 5365.71677977978u,1.5 5365.71777977978u,0 5376.46972022022u,0 5376.47072022022u,1.5 5377.447260260261u,1.5 5377.448260260261u,0 5378.4248003003u,0 5378.425800300301u,1.5 5380.37988038038u,1.5 5380.38088038038u,0 5381.357420420421u,0 5381.358420420421u,1.5 5392.110360860861u,1.5 5392.111360860861u,0 5393.0879009009u,0 5393.088900900901u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5411.661161661662u,0 5411.662161661662u,1.5 5412.638701701701u,1.5 5412.639701701702u,0 5415.571321821822u,0 5415.572321821822u,1.5 5417.526401901901u,1.5 5417.527401901902u,0 5418.503941941942u,0 5418.504941941942u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5434.144582582582u,0 5434.145582582582u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5442.942442942943u,0 5442.943442942943u,1.5 5443.919982982983u,1.5 5443.920982982983u,0 5457.605543543543u,0 5457.606543543543u,1.5 5458.583083583583u,1.5 5458.584083583583u,0 5460.538163663664u,0 5460.539163663664u,1.5 5461.515703703703u,1.5 5461.516703703704u,0 5466.403403903903u,0 5466.404403903904u,1.5 5467.380943943944u,1.5 5467.381943943944u,0 5468.358483983984u,0 5468.359483983984u,1.5 5469.336024024024u,1.5 5469.337024024024u,0 5471.291104104104u,0 5471.2921041041045u,1.5 5473.246184184184u,1.5 5473.247184184184u,0 5474.223724224224u,0 5474.224724224224u,1.5 5475.201264264265u,1.5 5475.202264264265u,0 5476.178804304304u,0 5476.1798043043045u,1.5 5478.133884384384u,1.5 5478.134884384384u,0 5479.1114244244245u,0 5479.112424424425u,1.5 5481.066504504504u,1.5 5481.0675045045045u,0 5482.044044544544u,0 5482.045044544544u,1.5 5490.841904904904u,1.5 5490.842904904905u,0 5491.819444944945u,0 5491.820444944945u,1.5 5493.774525025025u,1.5 5493.775525025025u,0 5494.752065065065u,0 5494.753065065065u,1.5 5497.684685185185u,1.5 5497.685685185185u,0 5498.662225225225u,0 5498.663225225225u,1.5 5511.370245745745u,1.5 5511.371245745745u,0 5512.347785785786u,0 5512.348785785786u,1.5 5520.168106106106u,1.5 5520.1691061061065u,0 5521.145646146146u,0 5521.146646146146u,1.5 5524.078266266267u,1.5 5524.079266266267u,0 5525.055806306306u,0 5525.0568063063065u,1.5 5527.9884264264265u,1.5 5527.989426426427u,0 5528.965966466467u,0 5528.966966466467u,1.5 5529.943506506506u,1.5 5529.9445065065065u,0 5533.853666666667u,0 5533.854666666667u,1.5 5534.831206706706u,1.5 5534.8322067067065u,0 5540.696446946947u,0 5540.697446946947u,1.5 5541.673986986987u,1.5 5541.674986986987u,0 5542.6515270270265u,0 5542.652527027027u,1.5 5543.629067067067u,1.5 5543.630067067067u,0 5557.3146276276275u,0 5557.315627627628u,1.5 5558.292167667668u,1.5 5558.293167667668u,0 5564.157407907907u,0 5564.1584079079075u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5569.045108108108u,0 5569.0461081081085u,1.5 5584.685748748749u,1.5 5584.686748748749u,0 5585.663288788789u,0 5585.664288788789u,1.5 5587.618368868869u,1.5 5587.619368868869u,0 5601.303929429429u,0 5601.30492942943u,1.5 5602.28146946947u,1.5 5602.28246946947u,0 5604.236549549549u,0 5604.237549549549u,1.5 5606.1916296296295u,1.5 5606.19262962963u,0 5607.16916966967u,0 5607.17016966967u,1.5 5616.94457007007u,1.5 5616.94557007007u,0 5617.92211011011u,0 5617.92311011011u,1.5 5619.87719019019u,1.5 5619.87819019019u,0 5620.8547302302295u,0 5620.85573023023u,1.5 5623.78735035035u,1.5 5623.78835035035u,0 5626.719970470471u,0 5626.720970470471u,1.5 5627.69751051051u,1.5 5627.6985105105105u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5648.225851351351u,1.5 5648.226851351351u,0 5650.180931431431u,0 5650.181931431432u,1.5 5652.136011511511u,1.5 5652.137011511511u,0 5659.956331831831u,0 5659.957331831832u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5662.888951951952u,0 5662.889951951952u,1.5 5673.641892392392u,1.5 5673.642892392392u,0 5674.619432432432u,0 5674.620432432433u,1.5 5675.596972472473u,1.5 5675.597972472473u,0 5685.372372872873u,0 5685.373372872873u,1.5 5686.349912912912u,1.5 5686.3509129129125u,0 5687.327452952953u,0 5687.328452952953u,1.5 5696.125313313313u,1.5 5696.126313313313u,0 5698.080393393393u,0 5698.081393393393u,1.5 5699.057933433433u,1.5 5699.058933433434u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5719.586274274275u,1.5 5719.587274274275u,0 5728.384134634634u,0 5728.385134634635u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5739.137075075075u,1.5 5739.138075075075u,0 5740.114615115115u,0 5740.115615115115u,1.5 5741.092155155155u,1.5 5741.093155155155u,0 5750.867555555555u,0 5750.868555555555u,1.5 5760.6429559559565u,1.5 5760.643955955957u,0 5762.598036036035u,0 5762.599036036036u,1.5 5763.575576076076u,1.5 5763.576576076076u,0 5769.440816316316u,0 5769.441816316316u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5780.1937567567575u,1.5 5780.194756756758u,0 5781.171296796797u,0 5781.172296796797u,1.5 5782.148836836836u,1.5 5782.149836836837u,0 5785.0814569569575u,0 5785.082456956958u,1.5 5786.058996996997u,1.5 5786.059996996997u,0 5791.924237237236u,0 5791.925237237237u,1.5 5794.8568573573575u,1.5 5794.857857357358u,0 5795.834397397397u,0 5795.835397397397u,1.5 5802.677177677678u,1.5 5802.678177677678u,0 5803.654717717717u,0 5803.655717717717u,1.5 5804.632257757758u,1.5 5804.633257757759u,0 5811.475038038037u,0 5811.476038038038u,1.5 5812.452578078078u,1.5 5812.453578078078u,0 5814.4076581581585u,0 5814.408658158159u,1.5 5816.362738238237u,1.5 5816.363738238238u,0 5817.340278278279u,0 5817.341278278279u,1.5 5827.115678678679u,1.5 5827.116678678679u,0 5833.958458958959u,0 5833.95945895896u,1.5 5834.935998998999u,1.5 5834.936998998999u,0 5836.891079079079u,0 5836.892079079079u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5839.823699199199u,0 5839.824699199199u,1.5 5849.5990995996u,1.5 5849.6000995996u,0 5850.576639639639u,0 5850.5776396396395u,1.5 5851.55417967968u,1.5 5851.55517967968u,0 5861.32958008008u,0 5861.33058008008u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5863.2846601601605u,0 5863.285660160161u,1.5 5864.2622002002u,1.5 5864.2632002002u,0 5865.239740240239u,0 5865.24074024024u,1.5 5866.217280280281u,1.5 5866.218280280281u,0 5867.19482032032u,0 5867.19582032032u,1.5 5877.947760760761u,1.5 5877.948760760762u,0 5878.925300800801u,0 5878.926300800801u,1.5 5879.90284084084u,1.5 5879.9038408408405u,0 5880.880380880881u,0 5880.881380880881u,1.5 5881.857920920921u,1.5 5881.858920920921u,0 5891.633321321321u,0 5891.634321321321u,1.5 5892.6108613613615u,1.5 5892.611861361362u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5896.521021521521u,1.5 5896.522021521521u,0 5897.4985615615615u,0 5897.499561561562u,1.5 5907.273961961962u,1.5 5907.274961961963u,0 5908.251502002002u,0 5908.252502002002u,1.5 5910.206582082082u,1.5 5910.207582082082u,0 5911.184122122122u,0 5911.185122122122u,1.5 5913.139202202202u,1.5 5913.140202202202u,0 5930.734922922923u,0 5930.735922922923u,1.5 5931.712462962963u,1.5 5931.713462962964u,0 5935.622623123123u,0 5935.623623123123u,1.5 5942.465403403403u,1.5 5942.466403403403u,0 5943.442943443443u,0 5943.4439434434435u,1.5 5962.993744244243u,1.5 5962.9947442442435u,0 5963.971284284285u,0 5963.972284284285u,1.5 5964.948824324324u,1.5 5964.949824324324u,0 5965.926364364364u,0 5965.927364364365u,1.5 5967.881444444444u,1.5 5967.882444444444u,0 5968.858984484485u,0 5968.859984484485u,1.5 5970.814064564564u,1.5 5970.815064564565u,0 5971.791604604605u,0 5971.792604604605u,1.5 5972.769144644644u,1.5 5972.7701446446445u,0 5973.746684684685u,0 5973.747684684685u,1.5 5974.724224724724u,1.5 5974.725224724724u,0 5976.679304804805u,0 5976.680304804805u,1.5 5977.656844844844u,1.5 5977.6578448448445u,0 5980.589464964965u,0 5980.590464964966u,1.5 5981.567005005005u,1.5 5981.568005005005u,0 5994.275025525525u,0 5994.276025525525u,1.5 5995.252565565565u,1.5 5995.253565565566u,0 6001.117805805806u,0 6001.118805805806u,1.5 6002.095345845845u,1.5 6002.0963458458455u,0 6013.825826326326u,0 6013.826826326326u,1.5 6014.803366366366u,1.5 6014.804366366367u,0 6019.691066566566u,0 6019.692066566567u,1.5 6020.668606606607u,1.5 6020.669606606607u,0 6024.578766766767u,0 6024.5797667667675u,1.5 6025.556306806807u,1.5 6025.557306806807u,0 6029.466466966967u,0 6029.467466966968u,1.5 6031.421547047046u,1.5 6031.4225470470465u,0 6033.376627127127u,0 6033.377627127127u,1.5 6034.354167167167u,1.5 6034.355167167168u,0 6035.331707207207u,0 6035.332707207207u,1.5 6037.286787287288u,1.5 6037.287787287288u,0 6038.264327327327u,0 6038.265327327327u,1.5 6061.7252882882885u,1.5 6061.726288288289u,0 6063.680368368368u,0 6063.681368368369u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6074.433308808809u,0 6074.434308808809u,1.5 6075.410848848848u,1.5 6075.411848848848u,0 6082.253629129129u,0 6082.254629129129u,1.5 6083.231169169169u,1.5 6083.2321691691695u,0 6084.208709209209u,0 6084.209709209209u,1.5 6085.186249249249u,1.5 6085.187249249249u,0 6087.141329329329u,0 6087.142329329329u,1.5 6088.118869369369u,1.5 6088.11986936937u,0 6090.073949449449u,0 6090.074949449449u,1.5 6091.0514894894895u,1.5 6091.05248948949u,0 6092.029029529529u,0 6092.030029529529u,1.5 6103.75951001001u,1.5 6103.76051001001u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6120.3776906906905u,0 6120.378690690691u,1.5 6121.35523073073u,1.5 6121.35623073073u,0 6122.332770770771u,0 6122.3337707707715u,1.5 6123.310310810811u,1.5 6123.311310810811u,0 6124.28785085085u,0 6124.28885085085u,1.5 6133.085711211211u,1.5 6133.086711211211u,0 6134.063251251251u,0 6134.064251251251u,1.5 6136.995871371371u,1.5 6136.9968713713715u,0 6147.748811811812u,0 6147.749811811812u,1.5 6148.726351851851u,1.5 6148.727351851851u,0 6149.7038918918915u,0 6149.704891891892u,1.5 6151.658971971972u,1.5 6151.6599719719725u,0 6152.636512012012u,0 6152.637512012012u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6161.434372372372u,0 6161.4353723723725u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6163.389452452452u,0 6163.390452452452u,1.5 6164.3669924924925u,1.5 6164.367992492493u,0 6172.187312812813u,0 6172.188312812813u,1.5 6173.164852852852u,1.5 6173.165852852852u,0 6175.119932932933u,0 6175.120932932933u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6195.648273773774u,0 6195.649273773774u,1.5 6196.625813813814u,1.5 6196.626813813814u,0 6197.603353853853u,0 6197.604353853853u,1.5 6207.378754254254u,1.5 6207.379754254254u,0 6217.154154654654u,0 6217.155154654654u,1.5 6219.109234734734u,1.5 6219.110234734734u,0 6220.086774774775u,0 6220.087774774775u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6230.839715215215u,0 6230.840715215215u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6238.660035535535u,0 6238.661035535535u,1.5 6239.637575575575u,1.5 6239.6385755755755u,0 6240.615115615616u,0 6240.616115615616u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6251.368056056055u,0 6251.369056056055u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6259.188376376376u,0 6259.1893763763765u,1.5 6260.165916416417u,1.5 6260.166916416417u,0 6261.143456456457u,0 6261.144456456457u,1.5 6262.120996496496u,1.5 6262.121996496497u,0 6263.098536536536u,0 6263.099536536536u,1.5 6267.0086966966965u,1.5 6267.009696696697u,0 6267.986236736736u,0 6267.987236736736u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6279.716717217217u,0 6279.717717217217u,1.5 6280.694257257258u,1.5 6280.695257257258u,0 6281.671797297297u,0 6281.672797297298u,1.5 6282.649337337337u,1.5 6282.650337337337u,0 6283.626877377377u,0 6283.627877377377u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6293.402277777778u,1.5 6293.403277777778u,0 6303.177678178178u,0 6303.178678178178u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6323.706019019019u,0 6323.707019019019u,1.5 6324.683559059059u,1.5 6324.684559059059u,0 6325.661099099099u,0 6325.6620990991u,1.5 6326.638639139139u,1.5 6326.639639139139u,0 6327.616179179179u,0 6327.617179179179u,1.5 6338.36911961962u,1.5 6338.37011961962u,0 6350.0996001001u,0 6350.100600100101u,1.5 6351.07714014014u,1.5 6351.07814014014u,0 6352.05468018018u,0 6352.05568018018u,1.5 6355.96484034034u,1.5 6355.96584034034u,0 6356.94238038038u,0 6356.94338038038u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6364.7627007007u,1.5 6364.763700700701u,0 6367.695320820821u,0 6367.696320820821u,1.5 6368.672860860861u,1.5 6368.673860860861u,0 6375.515641141141u,0 6375.516641141141u,1.5 6376.493181181181u,1.5 6376.494181181181u,0 6378.448261261262u,0 6378.449261261262u,1.5 6381.380881381381u,1.5 6381.381881381381u,0 6382.358421421422u,0 6382.359421421422u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6393.111361861862u,1.5 6393.112361861862u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6396.043981981982u,0 6396.044981981982u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6411.684622622623u,0 6411.685622622623u,1.5 6412.662162662663u,1.5 6412.663162662663u,0 6413.639702702702u,0 6413.640702702703u,1.5 6414.617242742742u,1.5 6414.618242742742u,0 6416.572322822823u,0 6416.573322822823u,1.5 6420.482482982983u,1.5 6420.483482982983u,0 6421.460023023023u,0 6421.461023023023u,1.5 6427.325263263264u,1.5 6427.326263263264u,0 6428.302803303303u,0 6428.3038033033035u,1.5 6432.212963463464u,1.5 6432.213963463464u,0 6433.190503503503u,0 6433.191503503504u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6436.1231236236235u,1.5 6436.124123623624u,0 6438.078203703703u,0 6438.079203703704u,1.5 6439.055743743743u,1.5 6439.056743743743u,0 6442.965903903903u,0 6442.966903903904u,1.5 6443.943443943944u,1.5 6443.944443943944u,0 6460.5616246246245u,0 6460.562624624625u,1.5 6461.539164664665u,1.5 6461.540164664665u,0 6466.426864864865u,0 6466.427864864865u,1.5 6467.404404904904u,1.5 6467.405404904905u,0 6468.381944944945u,0 6468.382944944945u,1.5 6469.359484984985u,1.5 6469.360484984985u,0 6470.337025025025u,0 6470.338025025025u,1.5 6471.314565065065u,1.5 6471.315565065065u,0 6472.292105105105u,0 6472.2931051051055u,1.5 6473.269645145145u,1.5 6473.270645145145u,0 6474.247185185185u,0 6474.248185185185u,1.5 6477.179805305305u,1.5 6477.1808053053055u,0 6478.157345345345u,0 6478.158345345345u,1.5 6483.045045545545u,1.5 6483.046045545545u,0 6484.022585585586u,0 6484.023585585586u,1.5 6485.0001256256255u,1.5 6485.001125625626u,0 6485.977665665666u,0 6485.978665665666u,1.5 6486.955205705705u,1.5 6486.9562057057055u,0 6487.932745745745u,0 6487.933745745745u,1.5 6489.8878258258255u,1.5 6489.888825825826u,0 6490.865365865866u,0 6490.866365865866u,1.5 6494.775526026026u,1.5 6494.776526026026u,0 6495.753066066066u,0 6495.754066066066u,1.5 6502.595846346346u,1.5 6502.596846346346u,0 6503.573386386386u,0 6503.574386386386u,1.5 6504.5509264264265u,1.5 6504.551926426427u,0 6505.528466466467u,0 6505.529466466467u,1.5 6509.4386266266265u,1.5 6509.439626626627u,0 6510.416166666667u,0 6510.417166666667u,1.5 6512.371246746747u,1.5 6512.372246746747u,0 6513.348786786787u,0 6513.349786786787u,1.5 6514.3263268268265u,1.5 6514.327326826827u,0 6515.303866866867u,0 6515.304866866867u,1.5 6516.281406906906u,1.5 6516.2824069069065u,0 6517.258946946947u,0 6517.259946946947u,1.5 6519.2140270270265u,1.5 6519.215027027027u,0 6520.191567067067u,0 6520.192567067067u,1.5 6521.169107107107u,1.5 6521.1701071071075u,0 6522.146647147147u,0 6522.147647147147u,1.5 6523.124187187187u,1.5 6523.125187187187u,0 6524.101727227227u,0 6524.102727227227u,1.5 6525.079267267268u,1.5 6525.080267267268u,0 6526.056807307307u,0 6526.0578073073075u,1.5 6528.011887387387u,1.5 6528.012887387387u,0 6529.966967467468u,0 6529.967967467468u,1.5 6531.922047547547u,1.5 6531.923047547547u,0 6532.899587587588u,0 6532.900587587588u,1.5 6533.8771276276275u,1.5 6533.878127627628u,0 6534.854667667668u,0 6534.855667667668u,1.5 6535.832207707707u,1.5 6535.8332077077075u,0 6538.7648278278275u,0 6538.765827827828u,1.5 6539.742367867868u,1.5 6539.743367867868u,0 6557.338088588589u,0 6557.339088588589u,1.5 6558.3156286286285u,1.5 6558.316628628629u,0 6560.270708708708u,0 6560.2717087087085u,1.5 6561.248248748749u,1.5 6561.249248748749u,0 6562.225788788789u,0 6562.226788788789u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6567.113488988989u,0 6567.114488988989u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.001189189189u,0 6572.002189189189u,1.5 6584.709209709709u,1.5 6584.7102097097095u,0 6585.68674974975u,0 6585.68774974975u,1.5 6586.66428978979u,1.5 6586.66528978979u,0 6588.61936986987u,0 6588.62036986987u,1.5 6591.55198998999u,1.5 6591.55298998999u,0 6602.30493043043u,0 6602.305930430431u,1.5 6603.282470470471u,1.5 6603.283470470471u,0 6606.215090590591u,0 6606.216090590591u,1.5 6608.170170670671u,1.5 6608.171170670671u,0 6609.14771071071u,0 6609.1487107107105u,1.5 6619.900651151151u,1.5 6619.901651151151u,0 6620.878191191191u,0 6620.879191191191u,1.5 6622.833271271272u,1.5 6622.834271271272u,0 6623.810811311311u,0 6623.811811311311u,1.5 6624.788351351351u,1.5 6624.789351351351u,0 6632.608671671672u,0 6632.609671671672u,1.5 6633.586211711711u,1.5 6633.5872117117115u,0 6634.563751751752u,0 6634.564751751752u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6640.428991991992u,1.5 6640.429991991992u,0 6641.4065320320315u,0 6641.407532032032u,1.5 6650.204392392392u,1.5 6650.205392392392u,0 6652.159472472473u,0 6652.160472472473u,1.5 6653.137012512512u,1.5 6653.138012512512u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6671.710273273274u,1.5 6671.711273273274u,0 6672.687813313313u,0 6672.688813313313u,1.5 6674.642893393393u,1.5 6674.643893393393u,0 6676.597973473474u,0 6676.598973473474u,1.5 6677.575513513513u,1.5 6677.576513513513u,0 6684.418293793794u,0 6684.419293793794u,1.5 6685.395833833833u,1.5 6685.396833833834u,0 6687.350913913913u,0 6687.351913913913u,1.5 6697.126314314314u,1.5 6697.127314314314u,0 6707.879254754755u,0 6707.880254754755u,1.5 6716.677115115115u,1.5 6716.678115115115u,0 6717.654655155155u,0 6717.655655155155u,1.5 6719.609735235234u,1.5 6719.610735235235u,0 6720.587275275276u,0 6720.588275275276u,1.5 6721.564815315315u,1.5 6721.565815315315u,0 6722.542355355355u,0 6722.543355355355u,1.5 6723.519895395395u,1.5 6723.520895395395u,0 6725.474975475476u,0 6725.475975475476u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6729.385135635635u,0 6729.386135635636u,1.5 6730.362675675676u,1.5 6730.363675675676u,0 6731.340215715715u,0 6731.341215715715u,1.5 6739.160536036035u,1.5 6739.161536036036u,0 6740.138076076076u,0 6740.139076076076u,1.5 6741.115616116116u,1.5 6741.116616116116u,0 6747.958396396396u,0 6747.959396396396u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5 6756.7562567567575u,1.5 6756.757256756758u,0 6757.733796796797u,0 6757.734796796797u,1.5 6758.711336836836u,1.5 6758.712336836837u,0 6759.688876876877u,0 6759.689876876877u,1.5 6762.621496996997u,1.5 6762.622496996997u,0 6770.441817317317u,0 6770.442817317317u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6780.217217717717u,1.5 6780.218217717717u,0 6792.925238238237u,0 6792.926238238238u,1.5 6802.700638638638u,1.5 6802.7016386386385u,0 6804.655718718718u,0 6804.656718718718u,1.5 6805.633258758759u,1.5 6805.63425875876u,0 6812.476039039038u,0 6812.477039039039u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6816.386199199199u,0 6816.387199199199u,1.5 6824.206519519519u,1.5 6824.207519519519u,0 6825.1840595595595u,0 6825.18505955956u,1.5 6826.1615995996u,1.5 6826.1625995996u,0 6827.139139639639u,0 6827.1401396396395u,1.5 6828.11667967968u,1.5 6828.11767967968u,0 6837.89208008008u,0 6837.89308008008u,1.5 6846.68994044044u,1.5 6846.6909404404405u,0 6847.667480480481u,0 6847.668480480481u,1.5 6850.600100600601u,1.5 6850.601100600601u,0 6854.510260760761u,0 6854.511260760762u,1.5 6855.487800800801u,1.5 6855.488800800801u,0 6864.285661161161u,0 6864.286661161162u,1.5 6865.263201201201u,1.5 6865.264201201201u,0 6866.24074124124u,0 6866.241741241241u,1.5 6873.083521521521u,1.5 6873.084521521521u,0 6874.0610615615615u,0 6874.062061561562u,1.5 6877.971221721721u,1.5 6877.972221721721u,0 6878.948761761762u,0 6878.949761761763u,1.5 6879.926301801802u,1.5 6879.927301801802u,0 6891.656782282283u,0 6891.657782282283u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5 6911.207583083083u,1.5 6911.208583083083u,0 6912.185123123123u,0 6912.186123123123u,1.5 6913.162663163163u,1.5 6913.163663163164u,0 6915.117743243242u,0 6915.1187432432425u,1.5 6916.095283283284u,1.5 6916.096283283284u,0 6929.780843843843u,0 6929.7818438438435u,1.5 6930.758383883884u,1.5 6930.759383883884u,0 6935.646084084084u,0 6935.647084084084u,1.5 6937.601164164164u,1.5 6937.602164164165u,0 6938.578704204204u,0 6938.579704204204u,1.5 6943.466404404404u,1.5 6943.467404404404u,0 6944.443944444444u,0 6944.444944444444u,1.5 6957.151964964965u,1.5 6957.152964964966u,0 6958.129505005005u,0 6958.130505005005u,1.5 6963.994745245244u,1.5 6963.9957452452445u,0 6964.972285285286u,0 6964.973285285286u,1.5 6965.949825325325u,1.5 6965.950825325325u,0 6966.927365365365u,0 6966.928365365366u,1.5 6968.882445445445u,1.5 6968.883445445445u,0 6971.815065565565u,0 6971.816065565566u,1.5 6972.792605605606u,1.5 6972.793605605606u,0 6973.770145645645u,0 6973.771145645645u,1.5 6974.747685685686u,1.5 6974.748685685686u,0 6975.725225725725u,0 6975.726225725725u,1.5 6976.702765765766u,1.5 6976.703765765767u,0 6980.612925925926u,0 6980.613925925926u,1.5 6981.590465965966u,1.5 6981.591465965967u,0 6986.478166166166u,0 6986.479166166167u,1.5 6987.455706206206u,1.5 6987.456706206206u,0 6988.433246246245u,0 6988.4342462462455u,1.5 6989.410786286287u,1.5 6989.411786286287u,0 6990.388326326326u,0 6990.389326326326u,1.5 6991.365866366366u,1.5 6991.366866366367u,0
vb23 b23 0 pwl 0,0  61.58452252252251u,0 61.58552252252252u,1.5 62.56206256256256u,1.5 62.563062562562564u,0 63.539602602602606u,0 63.54060260260261u,1.5 64.51714264264264u,1.5 64.51814264264264u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 67.44976276276276u,0 67.45076276276276u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 70.38238288288288u,1.5 70.38338288288288u,0 71.35992292292292u,0 71.36092292292292u,1.5 107.5289044044044u,1.5 107.5299044044044u,0 134.90002552552554u,0 134.9010255255255u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 137.83264564564567u,0 137.83364564564565u,1.5 163.2486866866867u,1.5 163.2496866866867u,0 184.7545675675676u,0 184.75556756756757u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 225.81124924924927u,0 225.81224924924925u,1.5 226.7887892892893u,1.5 226.78978928928927u,0 228.74386936936938u,0 228.74486936936935u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 271.75563113113117u,0 271.75663113113114u,1.5 291.3064319319319u,1.5 291.3074319319319u,0 292.28397197197194u,0 292.2849719719719u,1.5 294.23905205205205u,1.5 294.240052052052u,0 314.76739289289293u,0 314.7683928928929u,1.5 316.722472972973u,1.5 316.72347297297296u,0 317.700013013013u,0 317.701013013013u,1.5 334.31819369369373u,1.5 334.3191936936937u,0 335.2957337337337u,0 335.2967337337337u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 391.99305605605605u,1.5 391.994056056056u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 434.0272777777778u,0 434.02827777777776u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 436.9598978978979u,0 436.9608978978979u,1.5 442.82513813813813u,1.5 442.8261381381381u,0 443.80267817817816u,0 443.80367817817813u,1.5 447.7128383383383u,1.5 447.7138383383383u,0 448.69037837837834u,0 448.6913783783783u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 562.085023023023u,0 562.086023023023u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 567.9502632632633u,0 567.9512632632633u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 605.0967847847849u,0 605.0977847847848u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 608.0294049049048u,0 608.0304049049048u,1.5 633.445445945946u,1.5 633.4464459459459u,0 634.422985985986u,0 634.423985985986u,1.5 635.400526026026u,1.5 635.401526026026u,0 636.378066066066u,0 636.379066066066u,1.5 637.355606106106u,1.5 637.356606106106u,0 661.7941071071072u,0 661.7951071071071u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 665.7042672672673u,0 665.7052672672672u,1.5 684.277528028028u,1.5 684.278528028028u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 704.8058688688689u,0 704.8068688688688u,1.5 705.783408908909u,1.5 705.784408908909u,0 708.716029029029u,0 708.7170290290289u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 730.22190990991u,1.5 730.22290990991u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 791.8069324324325u,0 791.8079324324325u,1.5 813.3128133133133u,1.5 813.3138133133133u,0 815.2678933933934u,0 815.2688933933933u,1.5 816.2454334334335u,1.5 816.2464334334335u,0 817.2229734734735u,0 817.2239734734735u,1.5 818.2005135135136u,1.5 818.2015135135135u,0 834.8186941941941u,0 834.8196941941941u,1.5 835.7962342342342u,1.5 835.7972342342342u,0 836.7737742742743u,0 836.7747742742743u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 861.2122752752753u,1.5 861.2132752752752u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 866.0999754754755u,1.5 866.1009754754755u,0 895.4261766766766u,0 895.4271766766766u,1.5 929.6400780780781u,1.5 929.6410780780781u,0 930.6176181181181u,0 930.6186181181181u,1.5 934.5277782782782u,1.5 934.5287782782782u,0 935.5053183183182u,0 935.5063183183182u,1.5 936.4828583583584u,1.5 936.4838583583584u,0 939.4154784784785u,0 939.4164784784784u,1.5 940.3930185185185u,1.5 940.3940185185185u,0 1063.5630635635634u,0 1063.5640635635636u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1137.8561066066065u,0 1137.8571066066067u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1182.8229484484484u,0 1182.8239484484486u,1.5 1183.8004884884883u,1.5 1183.8014884884885u,0 1184.7780285285285u,0 1184.7790285285287u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1186.7331086086085u,0 1186.7341086086087u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1227.7897902902903u,0 1227.7907902902905u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1269.8240120120117u,1.5 1269.825012012012u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1289.3748128128127u,1.5 1289.375812812813u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1295.2400530530529u,1.5 1295.241053053053u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1336.2967347347346u,1.5 1336.2977347347348u,0 1337.2742747747748u,0 1337.275274774775u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1340.2068948948947u,0 1340.207894894895u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1363.6678558558558u,0 1363.668855855856u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1365.6229359359356u,0 1365.6239359359358u,1.5 1391.0389769769768u,1.5 1391.039976976977u,0 1392.016517017017u,0 1392.017517017017u,1.5 1392.9940570570568u,1.5 1392.995057057057u,0 1393.971597097097u,0 1393.9725970970972u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1395.926677177177u,0 1395.9276771771772u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1436.9833588588588u,0 1436.984358858859u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1440.8935190190189u,0 1440.894519019019u,1.5 1441.8710590590588u,1.5 1441.872059059059u,0 1442.848599099099u,0 1442.8495990990991u,1.5 1448.7138393393393u,1.5 1448.7148393393395u,0 1449.6913793793792u,0 1449.6923793793794u,1.5 1561.130943943944u,1.5 1561.1319439439442u,0 1562.108483983984u,0 1562.109483983984u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1566.018644144144u,0 1566.0196441441442u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1601.2100855855854u,0 1601.2110855855856u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1608.052865865866u,0 1608.053865865866u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1633.4689069069068u,1.5 1633.469906906907u,0 1634.446446946947u,0 1634.4474469469471u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1639.3341471471472u,0 1639.3351471471474u,1.5 1640.311687187187u,1.5 1640.3126871871873u,0 1658.884947947948u,0 1658.8859479479481u,1.5 1659.8624879879878u,1.5 1659.863487987988u,0 1663.7726481481482u,0 1663.7736481481484u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1686.256069069069u,0 1686.2570690690693u,1.5 1687.233609109109u,1.5 1687.2346091091092u,0 1706.7844099099098u,0 1706.78540990991u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1708.73948998999u,0 1708.7404899899902u,1.5 1711.67211011011u,1.5 1711.6731101101102u,0 1712.6496501501501u,0 1712.6506501501503u,1.5 1725.3576706706706u,1.5 1725.3586706706708u,0 1726.3352107107105u,0 1726.3362107107107u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1731.2229109109107u,0 1731.223910910911u,1.5 1732.2004509509509u,1.5 1732.201450950951u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1770.3245125125122u,1.5 1770.3255125125124u,0 1772.2795925925925u,0 1772.2805925925927u,1.5 1773.2571326326324u,1.5 1773.2581326326326u,0 1774.2346726726726u,0 1774.2356726726728u,1.5 1775.2122127127125u,1.5 1775.2132127127127u,0 1791.8303933933933u,0 1791.8313933933935u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1811.3811941941942u,1.5 1811.3821941941944u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1814.3138143143142u,0 1814.3148143143144u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1834.842155155155u,0 1834.8431551551553u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1861.235736236236u,1.5 1861.2367362362363u,0 1862.2132762762762u,0 1862.2142762762765u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1887.6293173173174u,0 1887.6303173173176u,1.5 1888.6068573573573u,1.5 1888.6078573573575u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1891.5394774774772u,1.5 1891.5404774774775u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1895.4496376376374u,0 1895.4506376376376u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1934.551239239239u,1.5 1934.5522392392393u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1939.4389394394395u,1.5 1939.4399394394397u,0 2058.698824324324u,0 2058.6998243243243u,1.5 2059.676364364364u,1.5 2059.677364364364u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2065.5416046046043u,1.5 2065.5426046046045u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2069.4517647647644u,0 2069.4527647647647u,1.5 2072.384384884885u,1.5 2072.3853848848853u,0 2073.3619249249246u,0 2073.3629249249248u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2107.575826326326u,0 2107.576826326326u,1.5 2108.553366366366u,1.5 2108.554366366366u,0 2112.463526526526u,0 2112.4645265265262u,1.5 2113.4410665665664u,1.5 2113.4420665665666u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2161.3405285285285u,1.5 2161.3415285285287u,0 2166.228228728729u,0 2166.229228728729u,1.5 2167.2057687687684u,1.5 2167.2067687687686u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2232.700951451451u,1.5 2232.7019514514514u,0 2233.6784914914915u,0 2233.6794914914917u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2271.802553053053u,1.5 2271.8035530530533u,0 2272.780093093093u,0 2272.781093093093u,1.5 2291.3533538538536u,1.5 2291.354353853854u,0 2292.330893893894u,0 2292.331893893894u,1.5 2294.285973973974u,1.5 2294.286973973974u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2317.746934934935u,1.5 2317.747934934935u,0 2318.724474974975u,0 2318.725474974975u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2361.736236736737u,1.5 2361.737236736737u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2365.646396896897u,0 2365.647396896897u,1.5 2388.1298178178176u,1.5 2388.130817817818u,0 2389.1073578578576u,0 2389.1083578578578u,1.5 2393.0175180180177u,1.5 2393.018518018018u,0 2393.995058058058u,0 2393.996058058058u,1.5 2394.972598098098u,1.5 2394.973598098098u,0 2395.9501381381383u,0 2395.9511381381385u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2398.882758258258u,0 2398.8837582582582u,1.5 2399.8602982982984u,1.5 2399.8612982982986u,0 2430.1640395395393u,0 2430.1650395395395u,1.5 2431.1415795795797u,1.5 2431.14257957958u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.0068198198196u,1.5 2437.00781981982u,0 2438.9618998999u,0 2438.9628998999u,1.5 2563.109484984985u,1.5 2563.1104849849853u,0 2564.0870250250246u,0 2564.0880250250248u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2571.907345345345u,1.5 2571.9083453453454u,0 2601.2335465465467u,0 2601.234546546547u,1.5 2602.2110865865866u,1.5 2602.212086586587u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2607.0987867867866u,0 2607.099786786787u,1.5 2636.424987987988u,1.5 2636.4259879879883u,0 2638.380068068068u,0 2638.381068068068u,1.5 2639.357608108108u,1.5 2639.358608108108u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2686.27953003003u,1.5 2686.28053003003u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2708.7629509509507u,1.5 2708.763950950951u,0 2709.740490990991u,0 2709.741490990991u,1.5 2726.3586716716713u,1.5 2726.3596716716715u,0 2727.3362117117117u,0 2727.337211711712u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2731.2463718718714u,1.5 2731.2473718718716u,0 2749.819632632633u,0 2749.820632632633u,1.5 2768.3928933933935u,1.5 2768.3938933933937u,0 2769.3704334334334u,0 2769.3714334334336u,1.5 2770.3479734734733u,1.5 2770.3489734734735u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2790.876314314314u,0 2790.8773143143144u,1.5 2791.853854354354u,1.5 2791.8548543543543u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2793.8089344344344u,1.5 2793.8099344344346u,0 2794.7864744744743u,0 2794.7874744744745u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2864.191817317317u,1.5 2864.1928173173173u,0 2889.607858358358u,0 2889.6088583583582u,1.5 2890.5853983983984u,1.5 2890.5863983983986u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2897.4281786786787u,1.5 2897.429178678679u,0 2898.4057187187186u,0 2898.406718718719u,1.5 2928.70945995996u,1.5 2928.71045995996u,0 2929.687u,0 2929.688u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2936.52978028028u,0 2936.5307802802804u,1.5 2937.50732032032u,1.5 2937.5083203203203u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2942.39502052052u,0 2942.3960205205203u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 3060.677365365365u,0 3060.678365365365u,1.5 3061.6549054054053u,1.5 3061.6559054054055u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3064.587525525525u,1.5 3064.5885255255253u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3069.4752257257255u,1.5 3069.4762257257257u,0 3070.4527657657654u,0 3070.4537657657656u,1.5 3074.3629259259255u,1.5 3074.3639259259257u,0 3075.340465965966u,0 3075.341465965966u,1.5 3098.8014269269265u,1.5 3098.8024269269267u,0 3099.778966966967u,0 3099.779966966967u,1.5 3102.711587087087u,1.5 3102.7125870870873u,0 3103.689127127127u,0 3103.690127127127u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3108.576827327327u,0 3108.577827327327u,1.5 3109.554367367367u,1.5 3109.555367367367u,0 3132.037788288288u,0 3132.0387882882883u,1.5 3133.0153283283285u,1.5 3133.0163283283287u,0 3134.9704084084083u,0 3134.9714084084085u,1.5 3136.9254884884886u,1.5 3136.9264884884888u,0 3137.9030285285285u,0 3137.9040285285287u,1.5 3161.3639894894895u,1.5 3161.3649894894897u,0 3162.3415295295295u,0 3162.3425295295297u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3164.2966096096093u,0 3164.2976096096095u,1.5 3165.2741496496496u,1.5 3165.27514964965u,0 3183.8474104104102u,0 3183.8484104104105u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3187.7575705705704u,0 3187.7585705705706u,1.5 3209.263451451451u,1.5 3209.2644514514514u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3269.870933933934u,0 3269.871933933934u,1.5 3270.848473973974u,1.5 3270.849473973974u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3273.781094094094u,0 3273.782094094094u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3312.8826956956955u,0 3312.8836956956957u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3315.8153158158157u,0 3315.816315815816u,1.5 3317.770395895896u,1.5 3317.771395895896u,0 3318.747935935936u,0 3318.748935935936u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3337.3211966966965u,0 3337.3221966966967u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3361.7596976976974u,0 3361.7606976976977u,1.5 3363.7147777777773u,1.5 3363.7157777777775u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3388.1532787787787u,1.5 3388.154278778779u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.0185190190186u,0 3394.019519019019u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3398.906219219219u,0 3398.9072192192193u,1.5 3399.883759259259u,1.5 3399.884759259259u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3437.0302807807807u,0 3437.031280780781u,1.5 3438.0078208208206u,1.5 3438.008820820821u,0 3438.9853608608605u,0 3438.9863608608607u,1.5 3561.1778658658654u,1.5 3561.1788658658656u,0 3562.155405905906u,0 3562.156405905906u,1.5 3564.110485985986u,1.5 3564.1114859859863u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.998186186186u,0 3568.9991861861863u,1.5 3569.975726226226u,1.5 3569.976726226226u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3609.0773278278275u,0 3609.0783278278277u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3681.4152907907906u,1.5 3681.4162907907908u,0 3682.392830830831u,0 3682.393830830831u,1.5 3685.3254509509507u,1.5 3685.326450950951u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3704.8762517517516u,0 3704.877251751752u,1.5 3705.8537917917915u,1.5 3705.8547917917917u,0 3707.8088718718714u,0 3707.8098718718716u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3728.3372127127127u,1.5 3728.338212712713u,0 3729.3147527527526u,0 3729.315752752753u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3733.2249129129127u,0 3733.225912912913u,1.5 3734.2024529529526u,1.5 3734.203452952953u,0 3746.9104734734733u,0 3746.9114734734735u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3770.3714344344344u,1.5 3770.3724344344346u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3862.260198198198u,1.5 3862.261198198198u,0 3864.2152782782778u,0 3864.216278278278u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3889.631319319319u,0 3889.6323193193193u,1.5 3890.608859359359u,1.5 3890.6098593593592u,0 3892.5639394394393u,0 3892.5649394394395u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 3929.710460960961u,1.5 3929.711460960961u,0 3930.688001001001u,0 3930.689001001001u,1.5 3931.665541041041u,1.5 3931.666541041041u,0 3932.643081081081u,0 3932.6440810810814u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3937.530781281281u,1.5 3937.5317812812814u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4069.4986866866866u,0 4069.499686686687u,1.5 4070.4762267267265u,1.5 4070.4772267267267u,0 4071.453766766767u,0 4071.454766766767u,1.5 4103.7125880880885u,1.5 4103.713588088089u,0 4104.690128128128u,0 4104.691128128128u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4131.083709209209u,0 4131.084709209209u,1.5 4132.061249249249u,1.5 4132.062249249249u,0 4136.948949449449u,0 4136.949949449449u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4139.881569569569u,0 4139.88256956957u,1.5 4160.40991041041u,1.5 4160.41091041041u,0 4161.38745045045u,0 4161.38845045045u,1.5 4162.3649904904905u,1.5 4162.365990490491u,0 4164.32007057057u,0 4164.321070570571u,1.5 4165.297610610611u,1.5 4165.298610610611u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4187.781031531531u,0 4187.782031531531u,1.5 4206.3542922922925u,1.5 4206.355292292293u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4210.264452452452u,0 4210.265452452452u,1.5 4211.2419924924925u,1.5 4211.242992492493u,0 4228.837713213213u,0 4228.838713213213u,1.5 4230.7927932932935u,1.5 4230.793793293294u,0 4231.770333333333u,0 4231.771333333333u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4266.961774774775u,0 4266.962774774775u,1.5 4267.939314814815u,1.5 4267.940314814815u,0 4271.849474974975u,0 4271.850474974975u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4315.838776776777u,0 4315.839776776777u,1.5 4316.816316816817u,1.5 4316.817316816817u,0 4317.793856856857u,0 4317.794856856857u,1.5 4334.412037537537u,1.5 4334.413037537537u,0 4335.389577577577u,0 4335.3905775775775u,1.5 4338.322197697697u,1.5 4338.323197697698u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4360.805618618619u,0 4360.806618618619u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4392.086899899899u,1.5 4392.0878998999u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.01952002002u,0 4395.02052002002u,1.5 4396.9746001001u,1.5 4396.975600100101u,0 4430.210961461462u,0 4430.211961461462u,1.5 4431.188501501501u,1.5 4431.189501501502u,0 4432.166041541541u,0 4432.167041541541u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4439.008821821822u,1.5 4439.009821821822u,0 4439.986361861862u,0 4439.987361861862u,1.5 4440.963901901901u,1.5 4440.964901901902u,0 4441.941441941942u,0 4441.942441941942u,1.5 4562.178866866867u,1.5 4562.179866866867u,0 4563.156406906906u,0 4563.1574069069065u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4569.021647147147u,0 4569.022647147147u,1.5 4569.999187187187u,1.5 4570.000187187187u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4607.145708708708u,1.5 4607.1467087087085u,0 4608.123248748749u,0 4608.124248748749u,1.5 4634.5168298298295u,1.5 4634.51782982983u,0 4635.49436986987u,0 4635.49536986987u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4640.38207007007u,0 4640.38307007007u,1.5 4641.35961011011u,1.5 4641.36061011011u,0 4659.932870870871u,0 4659.933870870871u,1.5 4660.91041091091u,1.5 4660.9114109109105u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4666.775651151151u,1.5 4666.776651151151u,0 4667.753191191191u,0 4667.754191191191u,1.5 4685.348911911911u,1.5 4685.3499119119115u,0 4686.326451951952u,0 4686.327451951952u,1.5 4687.303991991992u,1.5 4687.304991991992u,0 4688.2815320320315u,0 4688.282532032032u,1.5 4689.259072072072u,1.5 4689.260072072072u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4709.787412912912u,0 4709.7884129129125u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 4770.394895395395u,1.5 4770.395895395395u,0 4772.349975475476u,0 4772.350975475476u,1.5 4773.327515515515u,1.5 4773.328515515515u,0 4792.878316316316u,0 4792.879316316316u,1.5 4795.810936436436u,1.5 4795.811936436437u,0 4796.788476476477u,0 4796.789476476477u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4816.339277277278u,0 4816.340277277278u,1.5 4817.316817317317u,1.5 4817.317817317317u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4865.21627927928u,1.5 4865.21727927928u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4895.52002052052u,1.5 4895.52102052052u,0 4896.4975605605605u,0 4896.498560560561u,1.5 4930.711461961962u,1.5 4930.712461961963u,0 4931.689002002002u,0 4931.690002002002u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4935.599162162162u,1.5 4935.600162162163u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4939.509322322322u,0 4939.510322322322u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 5055.8365870870875u,0 5055.837587087088u,1.5 5056.814127127127u,1.5 5056.815127127127u,0 5059.746747247247u,0 5059.747747247247u,1.5 5060.724287287288u,1.5 5060.725287287288u,0 5061.701827327327u,0 5061.702827327327u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5067.567067567567u,1.5 5067.568067567568u,0 5068.544607607608u,0 5068.545607607608u,1.5 5071.477227727727u,1.5 5071.478227727727u,0 5072.454767767768u,0 5072.4557677677685u,1.5 5103.736049049048u,1.5 5103.737049049048u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5108.623749249249u,1.5 5108.624749249249u,0 5134.0397902902905u,0 5134.040790290291u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5136.97241041041u,0 5136.97341041041u,1.5 5137.94995045045u,1.5 5137.95095045045u,0 5138.9274904904905u,0 5138.928490490491u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5163.3659914914915u,0 5163.366991491492u,1.5 5164.343531531531u,1.5 5164.344531531531u,0 5181.939252252252u,0 5181.940252252252u,1.5 5182.9167922922925u,1.5 5182.917792292293u,0 5185.849412412412u,0 5185.850412412412u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5187.8044924924925u,0 5187.805492492493u,1.5 5207.3552932932935u,1.5 5207.356293293294u,0 5208.332833333333u,0 5208.333833333333u,1.5 5209.310373373373u,1.5 5209.3113733733735u,0 5210.287913413413u,0 5210.288913413413u,1.5 5211.265453453453u,1.5 5211.266453453453u,0 5228.861174174174u,0 5228.8621741741745u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5271.872935935936u,0 5271.873935935936u,1.5 5274.805556056056u,1.5 5274.806556056056u,0 5275.783096096096u,0 5275.784096096097u,1.5 5287.513576576576u,1.5 5287.5145765765765u,0 5288.491116616617u,0 5288.492116616617u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5316.839777777778u,0 5316.840777777778u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5359.851539539539u,0 5359.852539539539u,1.5 5360.829079579579u,1.5 5360.830079579579u,0 5365.71677977978u,0 5365.71777977978u,1.5 5392.110360860861u,1.5 5392.111360860861u,0 5393.0879009009u,0 5393.088900900901u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5433.167042542542u,0 5433.168042542542u,1.5 5434.144582582582u,1.5 5434.145582582582u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5442.942442942943u,1.5 5442.943442942943u,0 5443.919982982983u,0 5443.920982982983u,1.5 5557.3146276276275u,1.5 5557.315627627628u,0 5558.292167667668u,0 5558.293167667668u,1.5 5564.157407907907u,1.5 5564.1584079079075u,0 5568.067568068068u,0 5568.068568068068u,1.5 5569.045108108108u,1.5 5569.0461081081085u,0 5601.303929429429u,0 5601.30492942943u,1.5 5602.28146946947u,1.5 5602.28246946947u,0 5604.236549549549u,0 5604.237549549549u,1.5 5606.1916296296295u,1.5 5606.19262962963u,0 5607.16916966967u,0 5607.17016966967u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5659.956331831831u,0 5659.957331831832u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5662.888951951952u,0 5662.889951951952u,1.5 5685.372372872873u,1.5 5685.373372872873u,0 5686.349912912912u,0 5686.3509129129125u,1.5 5687.327452952953u,1.5 5687.328452952953u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5728.384134634634u,1.5 5728.385134634635u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5750.867555555555u,0 5750.868555555555u,1.5 5769.440816316316u,1.5 5769.441816316316u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5791.924237237236u,0 5791.925237237237u,1.5 5794.8568573573575u,1.5 5794.857857357358u,0 5795.834397397397u,0 5795.835397397397u,1.5 5811.475038038037u,1.5 5811.476038038038u,0 5812.452578078078u,0 5812.453578078078u,1.5 5814.4076581581585u,1.5 5814.408658158159u,0 5816.362738238237u,0 5816.363738238238u,1.5 5817.340278278279u,1.5 5817.341278278279u,0 5833.958458958959u,0 5833.95945895896u,1.5 5834.935998998999u,1.5 5834.936998998999u,0 5836.891079079079u,0 5836.892079079079u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5839.823699199199u,0 5839.824699199199u,1.5 5861.32958008008u,1.5 5861.33058008008u,0 5862.30712012012u,0 5862.30812012012u,1.5 5863.2846601601605u,1.5 5863.285660160161u,0 5864.2622002002u,0 5864.2632002002u,1.5 5865.239740240239u,1.5 5865.24074024024u,0 5866.217280280281u,0 5866.218280280281u,1.5 5867.19482032032u,1.5 5867.19582032032u,0 5891.633321321321u,0 5891.634321321321u,1.5 5892.6108613613615u,1.5 5892.611861361362u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5896.521021521521u,1.5 5896.522021521521u,0 5897.4985615615615u,0 5897.499561561562u,1.5 5930.734922922923u,1.5 5930.735922922923u,0 5931.712462962963u,0 5931.713462962964u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5942.465403403403u,0 5942.466403403403u,1.5 5943.442943443443u,1.5 5943.4439434434435u,0 6061.7252882882885u,0 6061.726288288289u,1.5 6063.680368368368u,1.5 6063.681368368369u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6074.433308808809u,1.5 6074.434308808809u,0 6075.410848848848u,0 6075.411848848848u,1.5 6103.75951001001u,1.5 6103.76051001001u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6133.085711211211u,0 6133.086711211211u,1.5 6134.063251251251u,1.5 6134.064251251251u,0 6136.995871371371u,0 6136.9968713713715u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6161.434372372372u,0 6161.4353723723725u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6163.389452452452u,0 6163.390452452452u,1.5 6164.3669924924925u,1.5 6164.367992492493u,0 6186.850413413413u,0 6186.851413413413u,1.5 6207.378754254254u,1.5 6207.379754254254u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6230.839715215215u,1.5 6230.840715215215u,0 6231.817255255255u,0 6231.818255255255u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6251.368056056055u,0 6251.369056056055u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6267.0086966966965u,0 6267.009696696697u,1.5 6267.986236736736u,1.5 6267.987236736736u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6293.402277777778u,1.5 6293.403277777778u,0 6315.885698698698u,0 6315.886698698699u,1.5 6338.36911961962u,1.5 6338.37011961962u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6364.7627007007u,0 6364.763700700701u,1.5 6367.695320820821u,1.5 6367.696320820821u,0 6368.672860860861u,0 6368.673860860861u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6393.111361861862u,1.5 6393.112361861862u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6396.043981981982u,0 6396.044981981982u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6427.325263263264u,0 6427.326263263264u,1.5 6428.302803303303u,1.5 6428.3038033033035u,0 6432.212963463464u,0 6432.213963463464u,1.5 6433.190503503503u,1.5 6433.191503503504u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6436.1231236236235u,0 6436.124123623624u,1.5 6438.078203703703u,1.5 6438.079203703704u,0 6439.055743743743u,0 6439.056743743743u,1.5 6442.965903903903u,1.5 6442.966903903904u,0 6443.943443943944u,0 6443.944443943944u,1.5 6557.338088588589u,1.5 6557.339088588589u,0 6558.3156286286285u,0 6558.316628628629u,1.5 6560.270708708708u,1.5 6560.2717087087085u,0 6561.248248748749u,0 6561.249248748749u,1.5 6562.225788788789u,1.5 6562.226788788789u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6566.135948948949u,0 6566.136948948949u,1.5 6567.113488988989u,1.5 6567.114488988989u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.001189189189u,1.5 6572.002189189189u,0 6602.30493043043u,0 6602.305930430431u,1.5 6603.282470470471u,1.5 6603.283470470471u,0 6606.215090590591u,0 6606.216090590591u,1.5 6608.170170670671u,1.5 6608.171170670671u,0 6609.14771071071u,0 6609.1487107107105u,1.5 6632.608671671672u,1.5 6632.609671671672u,0 6633.586211711711u,0 6633.5872117117115u,1.5 6634.563751751752u,1.5 6634.564751751752u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6640.428991991992u,0 6640.429991991992u,1.5 6641.4065320320315u,1.5 6641.407532032032u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6684.418293793794u,1.5 6684.419293793794u,0 6685.395833833833u,0 6685.396833833834u,1.5 6687.350913913913u,1.5 6687.351913913913u,0 6707.879254754755u,0 6707.880254754755u,1.5 6725.474975475476u,1.5 6725.475975475476u,0 6726.452515515515u,0 6726.453515515515u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6730.362675675676u,0 6730.363675675676u,1.5 6731.340215715715u,1.5 6731.341215715715u,0 6747.958396396396u,0 6747.959396396396u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5 6770.441817317317u,1.5 6770.442817317317u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6792.925238238237u,0 6792.926238238238u,1.5 6812.476039039038u,1.5 6812.477039039039u,0 6813.453579079079u,0 6813.454579079079u,1.5 6816.386199199199u,1.5 6816.387199199199u,0 6837.89208008008u,0 6837.89308008008u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6865.263201201201u,0 6865.264201201201u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6891.656782282283u,0 6891.657782282283u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5 6929.780843843843u,1.5 6929.7818438438435u,0 6930.758383883884u,0 6930.759383883884u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6937.601164164164u,0 6937.602164164165u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6943.466404404404u,0 6943.467404404404u,1.5 6944.443944444444u,1.5 6944.444944444444u,0
vb24 b24 0 pwl 0,0  107.5289044044044u,0 107.5299044044044u,1.5 163.2486866866867u,1.5 163.2496866866867u,0 208.21552852852852u,0 208.2165285285285u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 291.3064319319319u,0 291.3074319319319u,1.5 292.28397197197194u,1.5 292.2849719719719u,0 294.23905205205205u,0 294.240052052052u,1.5 334.31819369369373u,1.5 334.3191936936937u,0 335.2957337337337u,0 335.2967337337337u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 391.99305605605605u,0 391.994056056056u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 607.0518648648649u,0 607.0528648648649u,1.5 608.0294049049048u,1.5 608.0304049049048u,0 661.7941071071072u,0 661.7951071071071u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 665.7042672672673u,0 665.7052672672672u,1.5 704.8058688688689u,1.5 704.8068688688688u,0 705.783408908909u,0 705.784408908909u,1.5 708.716029029029u,1.5 708.7170290290289u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 791.8069324324325u,1.5 791.8079324324325u,0 834.8186941941941u,0 834.8196941941941u,1.5 835.7962342342342u,1.5 835.7972342342342u,0 836.7737742742743u,0 836.7747742742743u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 895.4261766766766u,1.5 895.4271766766766u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1289.3748128128127u,0 1289.375812812813u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1295.2400530530529u,0 1295.241053053053u,1.5 1336.2967347347346u,1.5 1336.2977347347348u,0 1337.2742747747748u,0 1337.275274774775u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1340.2068948948947u,0 1340.207894894895u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1391.0389769769768u,0 1391.039976976977u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1392.9940570570568u,0 1392.995057057057u,1.5 1393.971597097097u,1.5 1393.9725970970972u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1395.926677177177u,1.5 1395.9276771771772u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1601.2100855855854u,1.5 1601.2110855855856u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1608.052865865866u,1.5 1608.053865865866u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1658.884947947948u,0 1658.8859479479481u,1.5 1659.8624879879878u,1.5 1659.863487987988u,0 1663.7726481481482u,0 1663.7736481481484u,1.5 1706.7844099099098u,1.5 1706.78540990991u,0 1707.76194994995u,0 1707.76294994995u,1.5 1708.73948998999u,1.5 1708.7404899899902u,0 1711.67211011011u,0 1711.6731101101102u,1.5 1712.6496501501501u,1.5 1712.6506501501503u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1791.8303933933933u,1.5 1791.8313933933935u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1834.842155155155u,0 1834.8431551551553u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 1887.6293173173174u,1.5 1887.6303173173176u,0 1888.6068573573573u,0 1888.6078573573575u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1891.5394774774772u,0 1891.5404774774775u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1895.4496376376374u,1.5 1895.4506376376376u,0 2104.643206206206u,0 2104.644206206206u,1.5 2107.575826326326u,1.5 2107.576826326326u,0 2108.553366366366u,0 2108.554366366366u,1.5 2112.463526526526u,1.5 2112.4645265265262u,0 2113.4410665665664u,0 2113.4420665665666u,1.5 2161.3405285285285u,1.5 2161.3415285285287u,0 2166.228228728729u,0 2166.229228728729u,1.5 2167.2057687687684u,1.5 2167.2067687687686u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2291.3533538538536u,0 2291.354353853854u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2294.285973973974u,0 2294.286973973974u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2388.1298178178176u,0 2388.130817817818u,1.5 2389.1073578578576u,1.5 2389.1083578578578u,0 2393.0175180180177u,0 2393.018518018018u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2394.972598098098u,0 2394.973598098098u,1.5 2395.9501381381383u,1.5 2395.9511381381385u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2398.882758258258u,1.5 2398.8837582582582u,0 2399.8602982982984u,0 2399.8612982982986u,1.5 2601.2335465465467u,1.5 2601.234546546547u,0 2602.2110865865866u,0 2602.212086586587u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2607.0987867867866u,1.5 2607.099786786787u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2708.7629509509507u,0 2708.763950950951u,1.5 2709.740490990991u,1.5 2709.741490990991u,0 2749.819632632633u,0 2749.820632632633u,1.5 2790.876314314314u,1.5 2790.8773143143144u,0 2791.853854354354u,0 2791.8548543543543u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2793.8089344344344u,0 2793.8099344344346u,1.5 2794.7864744744743u,1.5 2794.7874744744745u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 2889.607858358358u,1.5 2889.6088583583582u,0 2890.5853983983984u,0 2890.5863983983986u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2897.4281786786787u,0 2897.429178678679u,1.5 2898.4057187187186u,1.5 2898.406718718719u,0 3098.8014269269265u,0 3098.8024269269267u,1.5 3099.778966966967u,1.5 3099.779966966967u,0 3102.711587087087u,0 3102.7125870870873u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3108.576827327327u,1.5 3108.577827327327u,0 3109.554367367367u,0 3109.555367367367u,1.5 3161.3639894894895u,1.5 3161.3649894894897u,0 3162.3415295295295u,0 3162.3425295295297u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3164.2966096096093u,0 3164.2976096096095u,1.5 3165.2741496496496u,1.5 3165.27514964965u,0 3209.263451451451u,0 3209.2644514514514u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3337.3211966966965u,0 3337.3221966966967u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3388.1532787787787u,0 3388.154278778779u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.0185190190186u,1.5 3394.019519019019u,0 3394.996059059059u,0 3394.997059059059u,1.5 3398.906219219219u,1.5 3398.9072192192193u,0 3399.883759259259u,0 3399.884759259259u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3609.0773278278275u,1.5 3609.0783278278277u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3704.8762517517516u,1.5 3704.877251751752u,0 3705.8537917917915u,0 3705.8547917917917u,1.5 3707.8088718718714u,1.5 3707.8098718718716u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3746.9104734734733u,0 3746.9114734734735u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 3889.631319319319u,1.5 3889.6323193193193u,0 3890.608859359359u,0 3890.6098593593592u,1.5 3892.5639394394393u,1.5 3892.5649394394395u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 4103.7125880880885u,0 4103.713588088089u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4106.645208208208u,0 4106.646208208208u,1.5 4160.40991041041u,1.5 4160.41091041041u,0 4161.38745045045u,0 4161.38845045045u,1.5 4162.3649904904905u,1.5 4162.365990490491u,0 4164.32007057057u,0 4164.321070570571u,1.5 4165.297610610611u,1.5 4165.298610610611u,0 4206.3542922922925u,0 4206.355292292293u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4210.264452452452u,1.5 4210.265452452452u,0 4211.2419924924925u,0 4211.242992492493u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4293.355355855856u,0 4293.356355855856u,1.5 4334.412037537537u,1.5 4334.413037537537u,0 4335.389577577577u,0 4335.3905775775775u,1.5 4338.322197697697u,1.5 4338.323197697698u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4392.086899899899u,0 4392.0878998999u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.01952002002u,1.5 4395.02052002002u,0 4396.9746001001u,0 4396.975600100101u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4607.145708708708u,0 4607.1467087087085u,1.5 4608.123248748749u,1.5 4608.124248748749u,0 4659.932870870871u,0 4659.933870870871u,1.5 4660.91041091091u,1.5 4660.9114109109105u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4666.775651151151u,1.5 4666.776651151151u,0 4667.753191191191u,0 4667.754191191191u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4709.787412912912u,1.5 4709.7884129129125u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 4792.878316316316u,1.5 4792.879316316316u,0 4795.810936436436u,0 4795.811936436437u,1.5 4796.788476476477u,1.5 4796.789476476477u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4895.52002052052u,0 4895.52102052052u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 5103.736049049048u,0 5103.737049049048u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5108.623749249249u,0 5108.624749249249u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5163.3659914914915u,0 5163.366991491492u,1.5 5164.343531531531u,1.5 5164.344531531531u,0 5207.3552932932935u,0 5207.356293293294u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5209.310373373373u,0 5209.3113733733735u,1.5 5210.287913413413u,1.5 5210.288913413413u,0 5211.265453453453u,0 5211.266453453453u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5287.513576576576u,0 5287.5145765765765u,1.5 5288.491116616617u,1.5 5288.492116616617u,0 5292.401276776777u,0 5292.402276776777u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5392.110360860861u,0 5392.111360860861u,1.5 5393.0879009009u,1.5 5393.088900900901u,0 5396.020521021021u,0 5396.021521021021u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5602.28146946947u,0 5602.28246946947u,1.5 5604.236549549549u,1.5 5604.237549549549u,0 5606.1916296296295u,0 5606.19262962963u,1.5 5607.16916966967u,1.5 5607.17016966967u,0 5659.956331831831u,0 5659.957331831832u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5662.888951951952u,0 5662.889951951952u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5750.867555555555u,0 5750.868555555555u,1.5 5791.924237237236u,1.5 5791.925237237237u,0 5794.8568573573575u,0 5794.857857357358u,1.5 5795.834397397397u,1.5 5795.835397397397u,0 5833.958458958959u,0 5833.95945895896u,1.5 5834.935998998999u,1.5 5834.936998998999u,0 5836.891079079079u,0 5836.892079079079u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5839.823699199199u,0 5839.824699199199u,1.5 5891.633321321321u,1.5 5891.634321321321u,0 5892.6108613613615u,0 5892.611861361362u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5896.521021521521u,0 5896.522021521521u,1.5 5897.4985615615615u,1.5 5897.499561561562u,0 6103.75951001001u,0 6103.76051001001u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6161.434372372372u,0 6161.4353723723725u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6163.389452452452u,0 6163.390452452452u,1.5 6164.3669924924925u,1.5 6164.367992492493u,0 6207.378754254254u,0 6207.379754254254u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6251.368056056055u,0 6251.369056056055u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6293.402277777778u,0 6293.403277777778u,1.5 6338.36911961962u,1.5 6338.37011961962u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6393.111361861862u,0 6393.112361861862u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6396.043981981982u,1.5 6396.044981981982u,0 6397.021522022022u,0 6397.022522022022u,1.5 6602.30493043043u,1.5 6602.305930430431u,0 6603.282470470471u,0 6603.283470470471u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6608.170170670671u,0 6608.171170670671u,1.5 6609.14771071071u,1.5 6609.1487107107105u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6747.958396396396u,0 6747.959396396396u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5 6792.925238238237u,1.5 6792.926238238238u,0 6837.89208008008u,0 6837.89308008008u,1.5 6891.656782282283u,1.5 6891.657782282283u,0 6892.634322322322u,0 6892.635322322322u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0
vb25 b25 0 pwl 0,0  163.2486866866867u,0 163.2496866866867u,1.5 249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 334.31819369369373u,0 334.3191936936937u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 337.2508138138138u,0 337.2518138138138u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 664.7267272272272u,0 664.7277272272272u,1.5 665.7042672672673u,1.5 665.7052672672672u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 834.8186941941941u,1.5 834.8196941941941u,0 835.7962342342342u,0 835.7972342342342u,1.5 836.7737742742743u,1.5 836.7747742742743u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1336.2967347347346u,0 1336.2977347347348u,1.5 1337.2742747747748u,1.5 1337.275274774775u,0 1338.251814814815u,0 1338.252814814815u,1.5 1340.2068948948947u,1.5 1340.207894894895u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1658.884947947948u,1.5 1658.8859479479481u,0 1659.8624879879878u,0 1659.863487987988u,1.5 1663.7726481481482u,1.5 1663.7736481481484u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 1834.842155155155u,1.5 1834.8431551551553u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 2161.3405285285285u,0 2161.3415285285287u,1.5 2166.228228728729u,1.5 2166.229228728729u,0 2167.2057687687684u,0 2167.2067687687686u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2749.819632632633u,0 2749.820632632633u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 3161.3639894894895u,0 3161.3649894894897u,1.5 3162.3415295295295u,1.5 3162.3425295295297u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3164.2966096096093u,1.5 3164.2976096096095u,0 3165.2741496496496u,0 3165.27514964965u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3337.3211966966965u,1.5 3337.3221966966967u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3746.9104734734733u,0 3746.9114734734735u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 4160.40991041041u,0 4160.41091041041u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4162.3649904904905u,0 4162.365990490491u,1.5 4164.32007057057u,1.5 4164.321070570571u,0 4165.297610610611u,0 4165.298610610611u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4334.412037537537u,0 4334.413037537537u,1.5 4335.389577577577u,1.5 4335.3905775775775u,0 4338.322197697697u,0 4338.323197697698u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4659.932870870871u,1.5 4659.933870870871u,0 4660.91041091091u,0 4660.9114109109105u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4666.775651151151u,0 4666.776651151151u,1.5 4667.753191191191u,1.5 4667.754191191191u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 5161.410911411411u,0 5161.411911411411u,1.5 5163.3659914914915u,1.5 5163.366991491492u,0 5164.343531531531u,0 5164.344531531531u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5339.323198698698u,0 5339.324198698699u,1.5 5659.956331831831u,1.5 5659.957331831832u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5662.888951951952u,1.5 5662.889951951952u,0 5750.867555555555u,0 5750.868555555555u,1.5 5833.958458958959u,1.5 5833.95945895896u,0 5834.935998998999u,0 5834.936998998999u,1.5 5836.891079079079u,1.5 5836.892079079079u,0 5837.868619119119u,0 5837.869619119119u,1.5 5839.823699199199u,1.5 5839.824699199199u,0 6160.456832332332u,0 6160.457832332332u,1.5 6161.434372372372u,1.5 6161.4353723723725u,0 6162.411912412412u,0 6162.412912412412u,1.5 6163.389452452452u,1.5 6163.390452452452u,0 6164.3669924924925u,0 6164.367992492493u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6251.368056056055u,0 6251.369056056055u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6338.36911961962u,0 6338.37011961962u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6747.958396396396u,0 6747.959396396396u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5 6837.89208008008u,1.5 6837.89308008008u,0
vb26 b26 0 pwl 0,0  249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 2250.296672172172u,0 2250.297672172172u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3746.9104734734733u,1.5 3746.9114734734735u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6251.368056056055u,1.5 6251.369056056055u,0 6252.345596096096u,0 6252.346596096097u,1.5 6747.958396396396u,1.5 6747.959396396396u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0

vbb21 bb21 0 pwl 0,0  2.93212012012012u,0 2.9331201201201202u,1.5 3.90966016016016u,1.5 3.9106601601601603u,0 10.75244044044044u,0 10.753440440440441u,1.5 11.72998048048048u,1.5 11.730980480480481u,0 17.59522072072072u,0 17.59622072072072u,1.5 18.572760760760765u,1.5 18.573760760760763u,0 21.50538088088088u,0 21.50638088088088u,1.5 22.482920920920925u,1.5 22.483920920920923u,0 27.370621121121122u,0 27.37162112112112u,1.5 28.348161161161162u,1.5 28.34916116116116u,0 29.325701201201202u,0 29.3267012012012u,1.5 30.303241241241246u,1.5 30.304241241241243u,0 32.25832132132132u,0 32.25932132132132u,1.5 37.146021521521526u,1.5 37.14702152152153u,0 38.12356156156156u,0 38.12456156156156u,1.5 40.07864164164164u,1.5 40.07964164164164u,0 41.05618168168168u,0 41.05718168168168u,1.5 42.03372172172172u,1.5 42.03472172172172u,0 43.01126176176176u,0 43.01226176176176u,1.5 46.92142192192192u,1.5 46.922421921921924u,0 47.89896196196196u,0 47.899961961961964u,1.5 49.85404204204204u,1.5 49.855042042042044u,0 51.80912212212212u,0 51.810122122122124u,1.5 52.786662162162166u,1.5 52.78766216216217u,0 56.69682232232232u,0 56.697822322322324u,1.5 57.67436236236236u,1.5 57.675362362362364u,0 61.58452252252251u,0 61.58552252252252u,1.5 62.56206256256256u,1.5 62.563062562562564u,0 63.539602602602606u,0 63.54060260260261u,1.5 64.51714264264264u,1.5 64.51814264264264u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 67.44976276276276u,0 67.45076276276276u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 70.38238288288288u,1.5 70.38338288288288u,0 71.35992292292292u,0 71.36092292292292u,1.5 73.315003003003u,1.5 73.316003003003u,0 75.27008308308308u,0 75.27108308308308u,1.5 77.22516316316316u,1.5 77.22616316316316u,0 78.2027032032032u,0 78.2037032032032u,1.5 79.18024324324324u,1.5 79.18124324324324u,0 81.13532332332332u,0 81.13632332332332u,1.5 83.0904034034034u,1.5 83.0914034034034u,0 85.04548348348348u,0 85.04648348348348u,1.5 86.02302352352352u,1.5 86.02402352352352u,0 88.95564364364364u,0 88.95664364364364u,1.5 89.9331836836837u,1.5 89.9341836836837u,0 90.91072372372372u,0 90.91172372372372u,1.5 92.8658038038038u,1.5 92.8668038038038u,0 93.84334384384384u,0 93.84434384384384u,1.5 96.77596396396396u,1.5 96.77696396396396u,0 107.5289044044044u,0 107.5299044044044u,1.5 114.37168468468468u,1.5 114.37268468468469u,0 115.34922472472472u,0 115.35022472472473u,1.5 116.32676476476476u,1.5 116.32776476476477u,0 120.23692492492492u,0 120.23792492492493u,1.5 121.21446496496498u,1.5 121.21546496496498u,0 122.19200500500502u,0 122.19300500500502u,1.5 124.14708508508508u,1.5 124.14808508508509u,0 125.12462512512512u,0 125.12562512512513u,1.5 129.0347852852853u,1.5 129.03578528528527u,0 130.01232532532532u,0 130.0133253253253u,1.5 130.98986536536538u,1.5 130.99086536536535u,0 134.90002552552554u,0 134.9010255255255u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 137.83264564564567u,0 137.83364564564565u,1.5 141.74280580580583u,1.5 141.7438058058058u,0 143.69788588588588u,0 143.69888588588586u,1.5 144.67542592592594u,1.5 144.6764259259259u,0 148.58558608608612u,0 148.5865860860861u,1.5 149.56312612612612u,1.5 149.5641261261261u,0 150.54066616616618u,0 150.54166616616615u,1.5 151.51820620620623u,1.5 151.5192062062062u,0 152.49574624624626u,0 152.49674624624623u,1.5 156.40590640640642u,1.5 156.4069064064064u,0 158.3609864864865u,0 158.36198648648647u,1.5 159.33852652652652u,1.5 159.3395265265265u,0 163.2486866866867u,0 163.2496866866867u,1.5 165.20376676676676u,1.5 165.20476676676674u,0 166.18130680680682u,0 166.1823068068068u,1.5 169.11392692692695u,1.5 169.11492692692693u,0 174.00162712712714u,0 174.0026271271271u,1.5 177.9117872872873u,1.5 177.91278728728727u,0 179.8668673673674u,0 179.86786736736738u,1.5 180.8444074074074u,1.5 180.84540740740738u,0 182.7994874874875u,0 182.8004874874875u,1.5 183.77702752752754u,1.5 183.7780275275275u,0 184.7545675675676u,0 184.75556756756757u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 190.6198078078078u,1.5 190.62080780780778u,0 192.57488788788788u,0 192.57588788788786u,1.5 193.55242792792794u,1.5 193.5534279279279u,0 194.529967967968u,0 194.53096796796797u,1.5 195.50750800800802u,1.5 195.508508008008u,0 197.4625880880881u,0 197.46358808808807u,1.5 201.37274824824826u,1.5 201.37374824824823u,0 203.32782832832834u,0 203.3288283283283u,1.5 204.3053683683684u,1.5 204.30636836836837u,0 208.21552852852852u,0 208.2165285285285u,1.5 215.05830880880882u,1.5 215.0593088088088u,0 217.0133888888889u,0 217.01438888888887u,1.5 217.99092892892892u,1.5 217.9919289289289u,0 218.96846896896898u,0 218.96946896896895u,1.5 221.90108908908908u,1.5 221.90208908908906u,0 223.85616916916916u,0 223.85716916916914u,1.5 224.83370920920922u,1.5 224.8347092092092u,0 225.81124924924927u,0 225.81224924924925u,1.5 226.7887892892893u,1.5 226.78978928928927u,0 228.74386936936938u,0 228.74486936936935u,1.5 234.60910960960962u,1.5 234.6101096096096u,0 239.4968098098098u,0 239.49780980980978u,1.5 242.42942992992997u,1.5 242.43042992992994u,0 243.40696996996996u,0 243.40796996996994u,1.5 245.36205005005007u,1.5 245.36305005005005u,0 247.31713013013015u,0 247.31813013013013u,1.5 248.29467017017018u,1.5 248.29567017017015u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 255.13745045045044u,1.5 255.13845045045042u,0 259.04761061061066u,0 259.04861061061064u,1.5 260.02515065065063u,1.5 260.0261506506506u,0 261.98023073073074u,0 261.9812307307307u,1.5 262.95777077077076u,1.5 262.95877077077074u,0 271.75563113113117u,0 271.75663113113114u,1.5 274.68825125125124u,1.5 274.6892512512512u,0 280.5534914914915u,0 280.5544914914915u,1.5 281.53103153153154u,1.5 281.5320315315315u,0 282.50857157157157u,0 282.50957157157154u,1.5 283.48611161161165u,1.5 283.4871116116116u,0 285.4411916916917u,0 285.4421916916917u,1.5 287.39627177177175u,1.5 287.3972717717717u,0 291.3064319319319u,0 291.3074319319319u,1.5 292.28397197197194u,1.5 292.2849719719719u,0 294.23905205205205u,0 294.240052052052u,1.5 299.12675225225223u,1.5 299.1277522522522u,0 302.0593723723724u,0 302.0603723723724u,1.5 303.03691241241245u,1.5 303.0379124124124u,0 304.9919924924925u,0 304.9929924924925u,1.5 305.9695325325325u,1.5 305.9705325325325u,0 306.9470725725726u,0 306.9480725725726u,1.5 308.90215265265266u,1.5 308.90315265265264u,0 314.76739289289293u,0 314.7683928928929u,1.5 316.722472972973u,1.5 316.72347297297296u,0 317.700013013013u,0 317.701013013013u,1.5 318.67755305305303u,1.5 318.678553053053u,0 319.6550930930931u,0 319.6560930930931u,1.5 320.63263313313314u,1.5 320.6336331331331u,0 325.5203333333333u,0 325.5213333333333u,1.5 326.4978733733734u,1.5 326.4988733733734u,0 327.47541341341343u,0 327.4764134134134u,1.5 329.4304934934935u,1.5 329.43149349349346u,0 331.3855735735736u,0 331.38657357357357u,1.5 332.3631136136136u,1.5 332.3641136136136u,0 333.3406536536537u,0 333.3416536536537u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 337.2508138138138u,0 337.2518138138138u,1.5 342.138514014014u,1.5 342.13951401401397u,0 343.1160540540541u,0 343.11705405405405u,1.5 345.0711341341341u,1.5 345.0721341341341u,0 346.0486741741742u,0 346.0496741741742u,1.5 347.02621421421424u,1.5 347.0272142142142u,0 348.9812942942943u,0 348.98229429429426u,1.5 349.9588343343343u,1.5 349.9598343343343u,0 350.9363743743744u,0 350.9373743743744u,1.5 351.9139144144144u,1.5 351.9149144144144u,0 352.8914544544545u,0 352.8924544544545u,1.5 353.8689944944945u,1.5 353.86999449449445u,0 354.8465345345345u,0 354.8475345345345u,1.5 355.8240745745746u,1.5 355.82507457457456u,0 357.7791546546547u,0 357.78015465465467u,1.5 358.7566946946947u,1.5 358.7576946946947u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 368.5320950950951u,1.5 368.53309509509506u,0 369.50963513513517u,0 369.51063513513515u,1.5 370.4871751751752u,1.5 370.4881751751752u,0 371.4647152152152u,0 371.4657152152152u,1.5 372.44225525525525u,1.5 372.4432552552552u,0 377.3299554554555u,0 377.33095545545547u,1.5 378.3074954954955u,1.5 378.3084954954955u,0 379.28503553553554u,0 379.2860355355355u,1.5 384.1727357357358u,1.5 384.17373573573576u,0 385.15027577577575u,0 385.15127577577573u,1.5 386.1278158158158u,1.5 386.12881581581576u,0 388.0828958958959u,0 388.08389589589586u,1.5 389.06043593593597u,1.5 389.06143593593595u,0 391.99305605605605u,0 391.994056056056u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 398.83583633633634u,1.5 398.8368363363363u,0 399.81337637637637u,0 399.81437637637634u,1.5 402.7459964964965u,1.5 402.7469964964965u,0 403.7235365365366u,0 403.72453653653656u,1.5 404.70107657657655u,1.5 404.70207657657653u,0 405.67861661661664u,0 405.6796166166166u,1.5 407.6336966966967u,1.5 407.63469669669666u,0 409.5887767767768u,0 409.5897767767768u,1.5 410.5663168168168u,1.5 410.5673168168168u,0 413.49893693693696u,0 413.49993693693693u,1.5 416.43155705705703u,1.5 416.432557057057u,0 417.40909709709706u,0 417.41009709709704u,1.5 418.38663713713714u,1.5 418.3876371371371u,0 419.36417717717717u,0 419.36517717717715u,1.5 421.3192572572573u,1.5 421.32025725725725u,0 422.29679729729736u,0 422.29779729729734u,1.5 423.27433733733733u,1.5 423.2753373373373u,0 424.25187737737735u,0 424.25287737737733u,1.5 426.20695745745746u,1.5 426.20795745745744u,0 427.18449749749755u,0 427.1854974974975u,1.5 428.16203753753757u,1.5 428.16303753753755u,0 433.04973773773776u,0 433.05073773773773u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 436.9598978978979u,0 436.9608978978979u,1.5 442.82513813813813u,1.5 442.8261381381381u,0 444.78021821821824u,0 444.7812182182182u,1.5 446.73529829829835u,1.5 446.7362982982983u,0 449.6679184184184u,0 449.6689184184184u,1.5 450.64545845845845u,1.5 450.6464584584584u,0 462.37593893893893u,0 462.3769389389389u,1.5 463.353478978979u,1.5 463.354478978979u,0 467.2636391391391u,0 467.2646391391391u,1.5 468.2411791791792u,1.5 468.2421791791792u,0 470.19625925925925u,0 470.1972592592592u,1.5 472.15133933933936u,1.5 472.15233933933933u,0 473.1288793793794u,0 473.12987937937936u,1.5 474.1064194194194u,1.5 474.1074194194194u,0 475.08395945945944u,0 475.0849594594594u,1.5 478.0165795795796u,1.5 478.0175795795796u,0 478.9941196196196u,0 478.9951196196196u,1.5 481.92673973973973u,1.5 481.9277397397397u,0 482.9042797797798u,0 482.9052797797798u,1.5 484.8593598598599u,1.5 484.8603598598599u,0 485.8368998998999u,0 485.83789989989987u,1.5 488.7695200200201u,1.5 488.77052002002006u,0 490.72460010010013u,0 490.7256001001001u,1.5 512.2304809809809u,1.5 512.2314809809809u,0 513.2080210210211u,0 513.209021021021u,1.5 514.1855610610611u,1.5 514.1865610610611u,0 517.1181811811812u,0 517.1191811811811u,1.5 518.0957212212213u,1.5 518.0967212212213u,0 519.0732612612613u,0 519.0742612612613u,1.5 520.0508013013012u,1.5 520.0518013013012u,0 521.0283413413413u,0 521.0293413413413u,1.5 525.9160415415415u,1.5 525.9170415415415u,0 526.8935815815815u,0 526.8945815815815u,1.5 527.8711216216217u,1.5 527.8721216216217u,0 529.8262017017017u,0 529.8272017017017u,1.5 531.7812817817818u,1.5 531.7822817817818u,0 534.7139019019019u,0 534.7149019019018u,1.5 535.6914419419419u,1.5 535.6924419419419u,0 537.646522022022u,0 537.647522022022u,1.5 538.6240620620621u,1.5 538.625062062062u,0 540.5791421421421u,0 540.5801421421421u,1.5 541.5566821821823u,1.5 541.5576821821822u,0 546.4443823823824u,0 546.4453823823824u,1.5 547.4219224224224u,1.5 547.4229224224224u,0 548.3994624624625u,0 548.4004624624624u,1.5 549.3770025025025u,1.5 549.3780025025025u,0 550.3545425425425u,0 550.3555425425425u,1.5 552.3096226226227u,1.5 552.3106226226226u,0 553.2871626626627u,0 553.2881626626627u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 562.085023023023u,0 562.086023023023u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 567.9502632632633u,0 567.9512632632633u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 570.8828833833834u,0 570.8838833833834u,1.5 571.8604234234234u,1.5 571.8614234234234u,0 573.8155035035035u,0 573.8165035035034u,1.5 574.7930435435435u,1.5 574.7940435435435u,0 577.7256636636637u,0 577.7266636636637u,1.5 579.6807437437437u,1.5 579.6817437437437u,0 580.6582837837839u,0 580.6592837837838u,1.5 587.501064064064u,1.5 587.502064064064u,0 588.4786041041041u,0 588.479604104104u,1.5 589.4561441441441u,1.5 589.4571441441441u,0 591.4112242242243u,0 591.4122242242242u,1.5 592.3887642642643u,1.5 592.3897642642643u,0 594.3438443443445u,0 594.3448443443444u,1.5 595.3213843843844u,1.5 595.3223843843843u,0 596.2989244244244u,0 596.2999244244244u,1.5 597.2764644644644u,1.5 597.2774644644644u,0 598.2540045045045u,0 598.2550045045044u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 607.0518648648649u,0 607.0528648648649u,1.5 608.0294049049048u,1.5 608.0304049049048u,0 610.962025025025u,0 610.963025025025u,1.5 611.939565065065u,1.5 611.940565065065u,0 613.8946451451452u,0 613.8956451451452u,1.5 614.8721851851852u,1.5 614.8731851851852u,0 615.8497252252253u,0 615.8507252252252u,1.5 619.7598853853854u,1.5 619.7608853853853u,0 620.7374254254254u,0 620.7384254254254u,1.5 621.7149654654654u,1.5 621.7159654654654u,0 622.6925055055054u,0 622.6935055055054u,1.5 623.6700455455456u,1.5 623.6710455455456u,0 626.6026656656657u,0 626.6036656656656u,1.5 627.5802057057057u,1.5 627.5812057057057u,0 629.5352857857858u,0 629.5362857857858u,1.5 633.445445945946u,1.5 633.4464459459459u,0 636.378066066066u,0 636.379066066066u,1.5 637.355606106106u,1.5 637.356606106106u,0 640.2882262262262u,0 640.2892262262262u,1.5 641.2657662662663u,1.5 641.2667662662662u,0 642.2433063063063u,0 642.2443063063063u,1.5 643.2208463463464u,1.5 643.2218463463464u,0 644.1983863863865u,0 644.1993863863864u,1.5 645.1759264264264u,1.5 645.1769264264263u,0 647.1310065065064u,0 647.1320065065064u,1.5 650.0636266266266u,1.5 650.0646266266266u,0 655.9288668668669u,0 655.9298668668669u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 664.7267272272272u,0 664.7277272272272u,1.5 665.7042672672673u,1.5 665.7052672672672u,0 668.6368873873874u,0 668.6378873873874u,1.5 672.5470475475475u,1.5 672.5480475475475u,0 674.5021276276276u,0 674.5031276276276u,1.5 675.4796676676676u,1.5 675.4806676676676u,0 678.4122877877878u,0 678.4132877877878u,1.5 680.3673678678679u,1.5 680.3683678678678u,0 681.344907907908u,0 681.345907907908u,1.5 682.3224479479479u,1.5 682.3234479479479u,0 683.299987987988u,0 683.3009879879879u,1.5 684.277528028028u,1.5 684.278528028028u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 689.1652282282282u,0 689.1662282282282u,1.5 690.1427682682682u,1.5 690.1437682682682u,0 691.1203083083084u,0 691.1213083083084u,1.5 693.0753883883884u,1.5 693.0763883883884u,0 694.0529284284285u,0 694.0539284284284u,1.5 696.9855485485485u,1.5 696.9865485485485u,0 697.9630885885886u,0 697.9640885885885u,1.5 698.9406286286286u,1.5 698.9416286286286u,0 701.8732487487488u,0 701.8742487487488u,1.5 703.8283288288288u,1.5 703.8293288288288u,0 705.783408908909u,0 705.784408908909u,1.5 709.693569069069u,1.5 709.694569069069u,0 713.6037292292292u,0 713.6047292292292u,1.5 715.5588093093094u,1.5 715.5598093093093u,0 716.5363493493494u,0 716.5373493493494u,1.5 718.4914294294294u,1.5 718.4924294294294u,0 719.4689694694696u,0 719.4699694694696u,1.5 720.4465095095095u,1.5 720.4475095095095u,0 723.3791296296296u,0 723.3801296296296u,1.5 725.3342097097097u,1.5 725.3352097097097u,0 726.3117497497498u,0 726.3127497497497u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 730.22190990991u,1.5 730.22290990991u,0 733.15453003003u,0 733.1555300300299u,1.5 734.1320700700701u,1.5 734.1330700700701u,0 736.0871501501501u,0 736.0881501501501u,1.5 739.0197702702703u,1.5 739.0207702702703u,0 743.9074704704706u,0 743.9084704704705u,1.5 745.8625505505505u,1.5 745.8635505505505u,0 746.8400905905905u,0 746.8410905905905u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 754.660410910911u,0 754.661410910911u,1.5 755.637950950951u,1.5 755.638950950951u,0 756.615490990991u,0 756.616490990991u,1.5 757.593031031031u,1.5 757.594031031031u,0 759.5481111111111u,0 759.5491111111111u,1.5 761.5031911911911u,1.5 761.5041911911911u,0 763.4582712712713u,0 763.4592712712713u,1.5 766.3908913913914u,1.5 766.3918913913914u,0 767.3684314314314u,0 767.3694314314314u,1.5 768.3459714714716u,1.5 768.3469714714715u,0 769.3235115115116u,0 769.3245115115116u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 774.2112117117117u,0 774.2122117117117u,1.5 775.1887517517517u,1.5 775.1897517517517u,0 776.1662917917918u,0 776.1672917917917u,1.5 778.1213718718719u,1.5 778.1223718718719u,0 779.098911911912u,0 779.0999119119119u,1.5 780.076451951952u,1.5 780.077451951952u,0 781.053991991992u,0 781.054991991992u,1.5 783.0090720720721u,1.5 783.010072072072u,0 785.9416921921921u,0 785.9426921921921u,1.5 786.9192322322323u,1.5 786.9202322322323u,0 787.8967722722723u,0 787.8977722722723u,1.5 791.8069324324325u,1.5 791.8079324324325u,0 796.6946326326326u,0 796.6956326326326u,1.5 797.6721726726727u,1.5 797.6731726726726u,0 798.6497127127127u,0 798.6507127127127u,1.5 799.6272527527527u,1.5 799.6282527527527u,0 800.6047927927928u,0 800.6057927927927u,1.5 801.5823328328329u,1.5 801.5833328328329u,0 802.5598728728729u,0 802.5608728728729u,1.5 803.5374129129129u,1.5 803.5384129129129u,0 804.514952952953u,0 804.515952952953u,1.5 806.4700330330331u,1.5 806.4710330330331u,0 808.4251131131131u,0 808.426113113113u,1.5 811.3577332332333u,1.5 811.3587332332332u,0 812.3352732732733u,0 812.3362732732733u,1.5 813.3128133133133u,1.5 813.3138133133133u,0 815.2678933933934u,0 815.2688933933933u,1.5 816.2454334334335u,1.5 816.2464334334335u,0 817.2229734734735u,0 817.2239734734735u,1.5 818.2005135135136u,1.5 818.2015135135135u,0 820.1555935935936u,0 820.1565935935936u,1.5 822.1106736736737u,1.5 822.1116736736736u,0 823.0882137137137u,0 823.0892137137137u,1.5 825.0432937937937u,1.5 825.0442937937937u,0 826.0208338338339u,0 826.0218338338339u,1.5 826.9983738738739u,1.5 826.9993738738739u,0 830.9085340340341u,0 830.9095340340341u,1.5 832.8636141141141u,1.5 832.864614114114u,0 833.8411541541541u,0 833.8421541541541u,1.5 834.8186941941941u,1.5 834.8196941941941u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 844.5940945945947u,0 844.5950945945947u,1.5 849.4817947947948u,1.5 849.4827947947948u,0 850.4593348348349u,0 850.4603348348348u,1.5 851.4368748748749u,1.5 851.4378748748749u,0 853.3919549549549u,0 853.3929549549549u,1.5 855.3470350350351u,1.5 855.3480350350351u,0 859.2571951951952u,0 859.2581951951952u,1.5 861.2122752752753u,1.5 861.2132752752752u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 866.0999754754755u,1.5 866.1009754754755u,0 869.0325955955957u,0 869.0335955955957u,1.5 871.9652157157157u,1.5 871.9662157157156u,0 872.9427557557557u,0 872.9437557557557u,1.5 873.9202957957958u,1.5 873.9212957957958u,0 875.8753758758759u,0 875.8763758758759u,1.5 877.8304559559559u,1.5 877.8314559559559u,0 878.8079959959961u,0 878.808995995996u,1.5 879.7855360360361u,1.5 879.7865360360361u,0 885.6507762762762u,0 885.6517762762762u,1.5 886.6283163163163u,1.5 886.6293163163162u,0 887.6058563563563u,0 887.6068563563563u,1.5 895.4261766766766u,1.5 895.4271766766766u,0 898.3587967967968u,0 898.3597967967968u,1.5 899.3363368368368u,1.5 899.3373368368368u,0 900.3138768768769u,0 900.3148768768768u,1.5 901.2914169169169u,1.5 901.2924169169169u,0 902.2689569569569u,0 902.2699569569569u,1.5 903.246496996997u,1.5 903.247496996997u,0 904.2240370370371u,0 904.225037037037u,1.5 905.2015770770771u,1.5 905.2025770770771u,0 907.1566571571572u,0 907.1576571571571u,1.5 910.0892772772772u,1.5 910.0902772772772u,0 913.9994374374375u,0 914.0004374374374u,1.5 915.9545175175175u,1.5 915.9555175175175u,0 918.8871376376377u,0 918.8881376376377u,1.5 919.8646776776777u,1.5 919.8656776776777u,0 920.8422177177176u,0 920.8432177177176u,1.5 921.8197577577578u,1.5 921.8207577577577u,0 922.7972977977978u,0 922.7982977977978u,1.5 928.6625380380381u,1.5 928.663538038038u,0 930.6176181181181u,0 930.6186181181181u,1.5 934.5277782782782u,1.5 934.5287782782782u,0 935.5053183183182u,0 935.5063183183182u,1.5 936.4828583583584u,1.5 936.4838583583584u,0 939.4154784784785u,0 939.4164784784784u,1.5 940.3930185185185u,1.5 940.3940185185185u,0 946.2582587587588u,0 946.2592587587587u,1.5 947.2357987987988u,1.5 947.2367987987988u,0 948.2133388388388u,0 948.2143388388388u,1.5 950.1684189189189u,1.5 950.1694189189188u,0 951.145958958959u,0 951.146958958959u,1.5 952.123498998999u,1.5 952.124498998999u,0 953.101039039039u,0 953.102039039039u,1.5 954.0785790790791u,1.5 954.079579079079u,0 955.0561191191191u,0 955.0571191191191u,1.5 960.9213593593594u,1.5 960.9223593593593u,0 962.8764394394394u,0 962.8774394394394u,1.5 964.8315195195195u,1.5 964.8325195195195u,0 965.8090595595596u,0 965.8100595595596u,1.5 968.7416796796797u,1.5 968.7426796796797u,0 970.6967597597597u,0 970.6977597597597u,1.5 972.6518398398398u,1.5 972.6528398398398u,0 973.6293798798798u,0 973.6303798798798u,1.5 974.60691991992u,1.5 974.6079199199199u,0 975.58445995996u,0 975.58545995996u,1.5 976.562u,1.5 976.563u,0 977.5395400400402u,0 977.5405400400401u,1.5 978.5170800800801u,1.5 978.51808008008u,0 982.4272402402403u,0 982.4282402402403u,1.5 983.4047802802802u,1.5 983.4057802802802u,0 984.3823203203203u,0 984.3833203203203u,1.5 985.3598603603602u,1.5 985.3608603603602u,0 986.3374004004004u,0 986.3384004004004u,1.5 987.3149404404405u,1.5 987.3159404404405u,0 988.2924804804804u,0 988.2934804804804u,1.5 989.2700205205206u,1.5 989.2710205205206u,0 993.1801806806807u,0 993.1811806806807u,1.5 994.1577207207208u,1.5 994.1587207207208u,0 997.0903408408409u,0 997.0913408408409u,1.5 998.0678808808808u,1.5 998.0688808808808u,0 999.045420920921u,0 999.0464209209209u,1.5 1001.9780410410411u,1.5 1001.9790410410411u,0 1011.7534414414415u,0 1011.7544414414415u,1.5 1014.6860615615615u,1.5 1014.6870615615614u,0 1021.5288418418419u,0 1021.5298418418419u,1.5 1022.5063818818818u,1.5 1022.5073818818818u,0 1023.4839219219219u,0 1023.4849219219219u,1.5 1025.4390020020019u,1.5 1025.440002002002u,0 1026.416542042042u,0 1026.4175420420422u,1.5 1027.394082082082u,1.5 1027.3950820820821u,0 1028.371622122122u,0 1028.3726221221223u,1.5 1029.349162162162u,1.5 1029.3501621621622u,0 1030.3267022022021u,0 1030.3277022022023u,1.5 1031.3042422422423u,1.5 1031.3052422422425u,0 1032.2817822822822u,0 1032.2827822822824u,1.5 1034.2368623623622u,1.5 1034.2378623623624u,0 1035.2144024024024u,0 1035.2154024024026u,1.5 1038.1470225225225u,1.5 1038.1480225225228u,0 1039.1245625625625u,0 1039.1255625625627u,1.5 1042.0571826826824u,1.5 1042.0581826826826u,0 1043.0347227227226u,0 1043.0357227227228u,1.5 1045.9673428428428u,1.5 1045.968342842843u,0 1046.9448828828827u,0 1046.9458828828829u,1.5 1047.9224229229228u,1.5 1047.923422922923u,0 1048.8999629629627u,0 1048.900962962963u,1.5 1049.8775030030029u,1.5 1049.878503003003u,0 1050.855043043043u,0 1050.8560430430432u,1.5 1051.832583083083u,1.5 1051.833583083083u,0 1052.810123123123u,0 1052.8111231231233u,1.5 1053.787663163163u,1.5 1053.7886631631632u,0 1055.7427432432432u,0 1055.7437432432434u,1.5 1056.7202832832832u,1.5 1056.7212832832834u,0 1063.5630635635634u,0 1063.5640635635636u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1073.338463963964u,1.5 1073.3394639639641u,0 1074.3160040040038u,0 1074.317004004004u,1.5 1077.248624124124u,1.5 1077.2496241241242u,0 1085.0689444444445u,0 1085.0699444444447u,1.5 1088.9791046046046u,1.5 1088.9801046046048u,0 1089.9566446446445u,0 1089.9576446446447u,1.5 1091.9117247247245u,1.5 1091.9127247247247u,0 1092.8892647647647u,0 1092.8902647647649u,1.5 1093.8668048048046u,1.5 1093.8678048048048u,0 1095.8218848848846u,0 1095.8228848848848u,1.5 1096.7994249249248u,1.5 1096.800424924925u,0 1099.732045045045u,0 1099.7330450450452u,1.5 1100.7095850850849u,1.5 1100.710585085085u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1112.4400655655656u,1.5 1112.4410655655659u,0 1113.4176056056056u,0 1113.4186056056058u,1.5 1115.3726856856854u,1.5 1115.3736856856856u,0 1120.2603858858856u,0 1120.2613858858858u,1.5 1121.2379259259258u,1.5 1121.238925925926u,0 1122.215465965966u,0 1122.216465965966u,1.5 1123.1930060060058u,1.5 1123.194006006006u,0 1124.170546046046u,0 1124.1715460460462u,1.5 1126.125626126126u,1.5 1126.1266261261262u,0 1128.080706206206u,0 1128.0817062062063u,1.5 1130.035786286286u,1.5 1130.0367862862863u,0 1131.0133263263263u,0 1131.0143263263265u,1.5 1131.9908663663664u,1.5 1131.9918663663666u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1137.8561066066065u,0 1137.8571066066067u,1.5 1140.7887267267265u,1.5 1140.7897267267267u,0 1141.7662667667666u,0 1141.7672667667669u,1.5 1143.7213468468467u,1.5 1143.722346846847u,0 1145.6764269269268u,0 1145.677426926927u,1.5 1146.653966966967u,1.5 1146.654966966967u,0 1148.609047047047u,0 1148.6100470470471u,1.5 1149.5865870870869u,1.5 1149.587587087087u,0 1150.564127127127u,0 1150.5651271271272u,1.5 1156.4293673673674u,1.5 1156.4303673673676u,0 1157.4069074074073u,0 1157.4079074074075u,1.5 1158.3844474474474u,1.5 1158.3854474474476u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1169.1373878878876u,1.5 1169.1383878878878u,0 1174.0250880880878u,0 1174.026088088088u,1.5 1175.9801681681681u,1.5 1175.9811681681683u,0 1176.957708208208u,0 1176.9587082082082u,1.5 1177.9352482482482u,1.5 1177.9362482482484u,0 1178.912788288288u,0 1178.9137882882883u,1.5 1179.8903283283282u,1.5 1179.8913283283284u,0 1180.8678683683684u,0 1180.8688683683686u,1.5 1183.8004884884883u,1.5 1183.8014884884885u,0 1184.7780285285285u,0 1184.7790285285287u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1186.7331086086085u,0 1186.7341086086087u,1.5 1191.6208088088085u,1.5 1191.6218088088087u,0 1193.5758888888888u,0 1193.576888888889u,1.5 1194.5534289289287u,1.5 1194.554428928929u,0 1195.5309689689689u,0 1195.531968968969u,1.5 1196.5085090090088u,1.5 1196.509509009009u,0 1197.486049049049u,0 1197.4870490490491u,1.5 1201.396209209209u,1.5 1201.3972092092092u,0 1202.3737492492492u,0 1202.3747492492494u,1.5 1203.3512892892893u,1.5 1203.3522892892895u,0 1204.3288293293292u,0 1204.3298293293294u,1.5 1205.3063693693693u,1.5 1205.3073693693696u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1212.1491496496496u,1.5 1212.1501496496498u,0 1213.1266896896898u,0 1213.12768968969u,1.5 1216.0593098098095u,1.5 1216.0603098098097u,0 1217.0368498498497u,0 1217.0378498498499u,1.5 1218.0143898898898u,1.5 1218.01538988989u,0 1218.9919299299297u,0 1218.99292992993u,1.5 1222.90209009009u,1.5 1222.9030900900902u,0 1223.87963013013u,0 1223.8806301301302u,1.5 1225.83471021021u,1.5 1225.8357102102102u,0 1227.7897902902903u,0 1227.7907902902905u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1234.6325705705706u,1.5 1234.6335705705708u,0 1239.5202707707706u,0 1239.5212707707708u,1.5 1241.4753508508506u,1.5 1241.4763508508508u,0 1242.4528908908908u,0 1242.453890890891u,1.5 1245.3855110110107u,1.5 1245.386511011011u,0 1247.340591091091u,0 1247.3415910910912u,1.5 1248.318131131131u,1.5 1248.3191311311311u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1256.1384514514514u,1.5 1256.1394514514516u,0 1259.0710715715716u,0 1259.0720715715718u,1.5 1261.0261516516516u,1.5 1261.0271516516518u,0 1262.0036916916918u,0 1262.004691691692u,1.5 1262.9812317317317u,1.5 1262.9822317317319u,0 1263.9587717717718u,0 1263.959771771772u,1.5 1264.9363118118117u,1.5 1264.937311811812u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1269.8240120120117u,1.5 1269.825012012012u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1274.711712212212u,1.5 1274.7127122122122u,0 1275.6892522522521u,0 1275.6902522522523u,1.5 1276.6667922922923u,1.5 1276.6677922922925u,0 1282.5320325325324u,0 1282.5330325325326u,1.5 1287.4197327327327u,1.5 1287.4207327327329u,0 1288.3972727727728u,0 1288.398272772773u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1296.217593093093u,0 1296.2185930930932u,1.5 1297.195133133133u,1.5 1297.1961331331331u,0 1298.172673173173u,0 1298.1736731731733u,1.5 1300.127753253253u,1.5 1300.1287532532533u,0 1301.1052932932932u,0 1301.1062932932934u,1.5 1302.0828333333332u,1.5 1302.0838333333334u,0 1303.0603733733733u,0 1303.0613733733735u,1.5 1305.0154534534533u,1.5 1305.0164534534536u,0 1306.9705335335334u,0 1306.9715335335336u,1.5 1308.9256136136135u,1.5 1308.9266136136137u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1320.656094094094u,1.5 1320.6570940940942u,0 1321.633634134134u,0 1321.634634134134u,1.5 1322.611174174174u,1.5 1322.6121741741742u,0 1324.566254254254u,0 1324.5672542542543u,1.5 1325.5437942942942u,1.5 1325.5447942942944u,0 1326.5213343343341u,0 1326.5223343343343u,1.5 1332.3865745745745u,1.5 1332.3875745745747u,0 1336.2967347347346u,0 1336.2977347347348u,1.5 1337.2742747747748u,1.5 1337.275274774775u,0 1338.251814814815u,0 1338.252814814815u,1.5 1340.2068948948947u,1.5 1340.207894894895u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1344.1170550550548u,1.5 1344.118055055055u,0 1345.094595095095u,0 1345.0955950950952u,1.5 1346.0721351351349u,1.5 1346.073135135135u,0 1350.9598353353351u,0 1350.9608353353353u,1.5 1352.9149154154154u,1.5 1352.9159154154156u,0 1353.8924554554553u,0 1353.8934554554555u,1.5 1354.8699954954955u,1.5 1354.8709954954957u,0 1355.8475355355354u,0 1355.8485355355356u,1.5 1356.8250755755755u,1.5 1356.8260755755757u,0 1358.7801556556556u,0 1358.7811556556558u,1.5 1359.7576956956957u,1.5 1359.758695695696u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1363.6678558558558u,0 1363.668855855856u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1365.6229359359356u,0 1365.6239359359358u,1.5 1370.5106361361359u,1.5 1370.511636136136u,0 1371.488176176176u,0 1371.4891761761762u,1.5 1372.4657162162162u,1.5 1372.4667162162164u,0 1378.3309564564563u,0 1378.3319564564565u,1.5 1380.2860365365364u,1.5 1380.2870365365366u,0 1381.2635765765765u,0 1381.2645765765767u,1.5 1383.2186566566565u,1.5 1383.2196566566568u,0 1384.1961966966967u,0 1384.197196696697u,1.5 1385.1737367367366u,1.5 1385.1747367367368u,0 1387.1288168168169u,0 1387.129816816817u,1.5 1388.1063568568568u,1.5 1388.107356856857u,0 1391.0389769769768u,0 1391.039976976977u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1392.9940570570568u,0 1392.995057057057u,1.5 1393.971597097097u,1.5 1393.9725970970972u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1395.926677177177u,1.5 1395.9276771771772u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1401.7919174174174u,1.5 1401.7929174174176u,0 1403.7469974974974u,0 1403.7479974974976u,1.5 1405.7020775775775u,1.5 1405.7030775775777u,0 1408.6346976976977u,0 1408.6356976976979u,1.5 1409.6122377377376u,1.5 1409.6132377377378u,0 1412.5448578578578u,0 1412.545857857858u,1.5 1413.522397897898u,1.5 1413.5233978978981u,0 1415.4774779779777u,0 1415.478477977978u,1.5 1416.4550180180179u,1.5 1416.456018018018u,0 1419.3876381381378u,0 1419.388638138138u,1.5 1420.365178178178u,1.5 1420.3661781781782u,0 1422.320258258258u,0 1422.3212582582582u,1.5 1423.2977982982982u,1.5 1423.2987982982984u,0 1424.275338338338u,0 1424.2763383383383u,1.5 1425.2528783783782u,1.5 1425.2538783783784u,0 1436.9833588588588u,0 1436.984358858859u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1440.8935190190189u,0 1440.894519019019u,1.5 1441.8710590590588u,1.5 1441.872059059059u,0 1443.826139139139u,0 1443.8271391391393u,1.5 1447.7362992992992u,1.5 1447.7372992992994u,0 1453.6015395395395u,0 1453.6025395395397u,1.5 1454.5790795795795u,1.5 1454.5800795795797u,0 1463.37693993994u,0 1463.3779399399402u,1.5 1464.35447997998u,1.5 1464.3554799799801u,0 1466.3095600600598u,0 1466.31056006006u,1.5 1467.2871001001u,1.5 1467.2881001001u,0 1468.26464014014u,0 1468.2656401401402u,1.5 1469.24218018018u,1.5 1469.2431801801802u,0 1476.0849604604603u,0 1476.0859604604605u,1.5 1478.0400405405405u,1.5 1478.0410405405407u,0 1479.0175805805804u,0 1479.0185805805806u,1.5 1482.9277407407408u,1.5 1482.928740740741u,0 1483.9052807807807u,0 1483.906280780781u,1.5 1486.8379009009009u,1.5 1486.838900900901u,0 1487.815440940941u,0 1487.8164409409412u,1.5 1488.792980980981u,1.5 1488.7939809809811u,0 1489.7705210210208u,0 1489.771521021021u,1.5 1493.680681181181u,1.5 1493.6816811811811u,0 1495.635761261261u,0 1495.6367612612612u,1.5 1496.6133013013011u,1.5 1496.6143013013013u,0 1498.5683813813812u,0 1498.5693813813814u,1.5 1499.5459214214213u,1.5 1499.5469214214215u,0 1500.5234614614612u,0 1500.5244614614614u,1.5 1501.5010015015014u,1.5 1501.5020015015016u,0 1502.4785415415415u,0 1502.4795415415417u,1.5 1506.3887017017016u,1.5 1506.3897017017018u,0 1508.3437817817817u,0 1508.3447817817819u,1.5 1512.253941941942u,1.5 1512.2549419419422u,0 1513.231481981982u,0 1513.2324819819821u,1.5 1514.209022022022u,1.5 1514.2100220220223u,0 1515.186562062062u,0 1515.1875620620622u,1.5 1521.0518023023021u,1.5 1521.0528023023023u,0 1522.0293423423423u,0 1522.0303423423425u,1.5 1525.9395025025024u,1.5 1525.9405025025026u,0 1528.8721226226226u,0 1528.8731226226228u,1.5 1529.8496626626625u,1.5 1529.8506626626627u,0 1530.8272027027026u,0 1530.8282027027028u,1.5 1531.8047427427427u,1.5 1531.805742742743u,0 1534.7373628628627u,0 1534.738362862863u,1.5 1535.7149029029028u,1.5 1535.715902902903u,0 1537.669982982983u,0 1537.670982982983u,1.5 1538.647523023023u,1.5 1538.6485230230232u,0 1539.625063063063u,0 1539.6260630630632u,1.5 1542.557683183183u,1.5 1542.5586831831831u,0 1546.4678433433432u,0 1546.4688433433435u,1.5 1547.4453833833832u,1.5 1547.4463833833834u,0 1549.4004634634632u,0 1549.4014634634634u,1.5 1550.3780035035034u,1.5 1550.3790035035036u,0 1551.3555435435435u,0 1551.3565435435437u,1.5 1552.3330835835834u,1.5 1552.3340835835836u,0 1553.3106236236235u,0 1553.3116236236237u,1.5 1556.2432437437437u,1.5 1556.244243743744u,0 1557.2207837837836u,0 1557.2217837837838u,1.5 1561.130943943944u,1.5 1561.1319439439442u,0 1563.086024024024u,0 1563.0870240240242u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1566.018644144144u,0 1566.0196441441442u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1577.7491246246245u,0 1577.7501246246247u,1.5 1581.6592847847846u,1.5 1581.6602847847848u,0 1582.6368248248248u,0 1582.637824824825u,1.5 1583.614364864865u,1.5 1583.6153648648651u,0 1584.5919049049048u,0 1584.592904904905u,1.5 1587.524525025025u,1.5 1587.5255250250252u,0 1589.479605105105u,0 1589.4806051051053u,1.5 1590.457145145145u,1.5 1590.4581451451452u,0 1596.3223853853851u,0 1596.3233853853853u,1.5 1598.2774654654654u,1.5 1598.2784654654656u,0 1599.2550055055053u,0 1599.2560055055055u,1.5 1600.2325455455455u,1.5 1600.2335455455457u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1610.9854859859859u,0 1610.986485985986u,1.5 1611.963026026026u,1.5 1611.9640260260262u,0 1612.9405660660661u,0 1612.9415660660663u,1.5 1614.8956461461462u,1.5 1614.8966461461464u,0 1615.8731861861859u,0 1615.874186186186u,1.5 1616.850726226226u,1.5 1616.8517262262262u,0 1617.8282662662662u,0 1617.8292662662664u,1.5 1619.7833463463462u,1.5 1619.7843463463464u,0 1620.7608863863861u,0 1620.7618863863863u,1.5 1621.7384264264263u,1.5 1621.7394264264265u,0 1622.7159664664664u,0 1622.7169664664666u,1.5 1623.6935065065063u,1.5 1623.6945065065065u,0 1624.6710465465464u,0 1624.6720465465467u,1.5 1625.6485865865864u,1.5 1625.6495865865866u,0 1628.5812067067066u,0 1628.5822067067068u,1.5 1629.5587467467467u,1.5 1629.559746746747u,0 1630.5362867867866u,0 1630.5372867867868u,1.5 1633.4689069069068u,1.5 1633.469906906907u,0 1634.446446946947u,0 1634.4474469469471u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1639.3341471471472u,0 1639.3351471471474u,1.5 1640.311687187187u,1.5 1640.3126871871873u,0 1642.2667672672671u,0 1642.2677672672673u,1.5 1644.2218473473472u,1.5 1644.2228473473474u,0 1645.199387387387u,0 1645.2003873873873u,1.5 1649.1095475475474u,1.5 1649.1105475475476u,0 1651.0646276276275u,0 1651.0656276276277u,1.5 1652.0421676676676u,1.5 1652.0431676676678u,0 1655.9523278278277u,0 1655.953327827828u,1.5 1656.9298678678679u,1.5 1656.930867867868u,0 1657.9074079079078u,0 1657.908407907908u,1.5 1658.884947947948u,1.5 1658.8859479479481u,0 1660.840028028028u,0 1660.8410280280282u,1.5 1664.750188188188u,1.5 1664.7511881881883u,0 1667.682808308308u,0 1667.6838083083082u,1.5 1674.5255885885883u,1.5 1674.5265885885885u,0 1680.3908288288287u,0 1680.391828828829u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1686.256069069069u,0 1686.2570690690693u,1.5 1687.233609109109u,1.5 1687.2346091091092u,0 1691.1437692692691u,0 1691.1447692692693u,1.5 1696.0314694694694u,1.5 1696.0324694694696u,0 1697.9865495495494u,0 1697.9875495495496u,1.5 1698.9640895895895u,1.5 1698.9650895895898u,0 1701.8967097097095u,0 1701.8977097097097u,1.5 1702.8742497497497u,1.5 1702.8752497497499u,0 1703.8517897897898u,0 1703.85278978979u,1.5 1704.8293298298297u,1.5 1704.83032982983u,0 1705.8068698698698u,0 1705.80786986987u,1.5 1706.7844099099098u,1.5 1706.78540990991u,0 1707.76194994995u,0 1707.76294994995u,1.5 1708.73948998999u,1.5 1708.7404899899902u,0 1710.69457007007u,0 1710.6955700700703u,1.5 1717.5373503503502u,1.5 1717.5383503503504u,0 1718.5148903903903u,0 1718.5158903903905u,1.5 1719.4924304304302u,1.5 1719.4934304304304u,0 1727.3127507507506u,0 1727.3137507507508u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1731.2229109109107u,0 1731.223910910911u,1.5 1732.2004509509509u,1.5 1732.201450950951u,0 1733.177990990991u,0 1733.1789909909912u,1.5 1739.0432312312312u,1.5 1739.0442312312314u,0 1740.0207712712713u,0 1740.0217712712715u,1.5 1740.998311311311u,1.5 1740.9993113113112u,0 1741.9758513513511u,0 1741.9768513513513u,1.5 1743.9309314314312u,1.5 1743.9319314314314u,0 1745.8860115115112u,0 1745.8870115115114u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1755.6614119119117u,0 1755.662411911912u,1.5 1760.549112112112u,1.5 1760.5501121121122u,0 1762.5041921921922u,0 1762.5051921921925u,1.5 1763.4817322322322u,1.5 1763.4827322322324u,0 1765.4368123123122u,0 1765.4378123123124u,1.5 1770.3245125125122u,1.5 1770.3255125125124u,0 1772.2795925925925u,0 1772.2805925925927u,1.5 1773.2571326326324u,1.5 1773.2581326326326u,0 1774.2346726726726u,0 1774.2356726726728u,1.5 1776.1897527527526u,1.5 1776.1907527527528u,0 1777.1672927927928u,0 1777.168292792793u,1.5 1778.1448328328327u,1.5 1778.1458328328329u,0 1779.1223728728728u,0 1779.123372872873u,1.5 1782.054992992993u,1.5 1782.0559929929932u,0 1787.9202332332331u,0 1787.9212332332334u,1.5 1788.8977732732733u,1.5 1788.8987732732735u,0 1789.8753133133132u,0 1789.8763133133134u,1.5 1791.8303933933933u,1.5 1791.8313933933935u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1797.6956336336334u,0 1797.6966336336336u,1.5 1798.6731736736735u,1.5 1798.6741736736737u,0 1799.6507137137135u,0 1799.6517137137137u,1.5 1800.6282537537536u,1.5 1800.6292537537538u,0 1801.6057937937937u,0 1801.606793793794u,1.5 1804.5384139139137u,1.5 1804.539413913914u,0 1806.493493993994u,0 1806.4944939939942u,1.5 1807.471034034034u,1.5 1807.472034034034u,0 1808.448574074074u,0 1808.4495740740742u,1.5 1809.426114114114u,1.5 1809.4271141141141u,0 1810.403654154154u,0 1810.4046541541543u,1.5 1811.3811941941942u,1.5 1811.3821941941944u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1814.3138143143142u,0 1814.3148143143144u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1820.1790545545543u,0 1820.1800545545545u,1.5 1821.1565945945945u,1.5 1821.1575945945947u,0 1822.1341346346344u,0 1822.1351346346346u,1.5 1823.1116746746745u,1.5 1823.1126746746747u,0 1824.0892147147147u,0 1824.0902147147149u,1.5 1826.0442947947947u,1.5 1826.045294794795u,0 1827.9993748748748u,0 1828.000374874875u,1.5 1829.9544549549548u,1.5 1829.955454954955u,0 1830.931994994995u,0 1830.9329949949952u,1.5 1831.9095350350349u,1.5 1831.910535035035u,0 1832.887075075075u,0 1832.8880750750752u,1.5 1833.8646151151152u,1.5 1833.8656151151154u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1843.6400155155154u,0 1843.6410155155156u,1.5 1844.6175555555553u,1.5 1844.6185555555555u,0 1845.5950955955955u,0 1845.5960955955957u,1.5 1851.4603358358356u,1.5 1851.4613358358358u,0 1855.370495995996u,0 1855.3714959959962u,1.5 1857.325576076076u,1.5 1857.3265760760762u,0 1858.3031161161161u,0 1858.3041161161163u,1.5 1859.280656156156u,1.5 1859.2816561561563u,0 1860.2581961961962u,0 1860.2591961961964u,1.5 1861.235736236236u,1.5 1861.2367362362363u,0 1862.2132762762762u,0 1862.2142762762765u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1867.1009764764763u,0 1867.1019764764765u,1.5 1868.0785165165164u,1.5 1868.0795165165166u,0 1871.0111366366364u,0 1871.0121366366366u,1.5 1872.9662167167166u,1.5 1872.9672167167168u,0 1873.9437567567566u,0 1873.9447567567568u,1.5 1876.8763768768767u,1.5 1876.877376876877u,0 1877.853916916917u,0 1877.854916916917u,1.5 1878.8314569569568u,1.5 1878.832456956957u,0 1880.7865370370369u,0 1880.787537037037u,1.5 1882.7416171171171u,1.5 1882.7426171171173u,0 1884.6966971971972u,0 1884.6976971971974u,1.5 1885.674237237237u,1.5 1885.6752372372373u,0 1888.6068573573573u,0 1888.6078573573575u,1.5 1889.5843973973974u,1.5 1889.5853973973976u,0 1891.5394774774772u,0 1891.5404774774775u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1895.4496376376374u,1.5 1895.4506376376376u,0 1900.3373378378376u,0 1900.3383378378378u,1.5 1901.3148778778777u,1.5 1901.315877877878u,0 1903.2699579579578u,0 1903.270957957958u,1.5 1906.202578078078u,1.5 1906.2035780780782u,0 1907.1801181181181u,0 1907.1811181181183u,1.5 1913.0453583583583u,1.5 1913.0463583583585u,0 1914.0228983983984u,0 1914.0238983983986u,1.5 1915.0004384384383u,1.5 1915.0014384384385u,0 1921.8432187187186u,0 1921.8442187187188u,1.5 1924.7758388388386u,1.5 1924.7768388388388u,0 1925.7533788788787u,0 1925.754378878879u,1.5 1928.685998998999u,1.5 1928.6869989989991u,0 1929.6635390390388u,0 1929.664539039039u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1934.551239239239u,1.5 1934.5522392392393u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1939.4389394394395u,1.5 1939.4399394394397u,0 1942.3715595595593u,0 1942.3725595595595u,1.5 1943.3490995995994u,1.5 1943.3500995995996u,0 1947.2592597597595u,0 1947.2602597597597u,1.5 1948.2367997997997u,1.5 1948.2377997997999u,0 1950.1918798798797u,0 1950.19287987988u,1.5 1951.1694199199198u,1.5 1951.17041991992u,0 1952.1469599599598u,0 1952.14795995996u,1.5 1953.1245u,1.5 1953.1255u,0 1954.10204004004u,0 1954.1030400400402u,1.5 1955.0795800800802u,1.5 1955.0805800800804u,0 1956.0571201201199u,0 1956.05812012012u,1.5 1959.9672802802804u,1.5 1959.9682802802806u,0 1961.9223603603602u,0 1961.9233603603604u,1.5 1967.7876006006004u,1.5 1967.7886006006006u,0 1969.7426806806807u,0 1969.7436806806809u,1.5 1970.7202207207204u,1.5 1970.7212207207206u,0 1971.6977607607605u,0 1971.6987607607607u,1.5 1972.6753008008006u,1.5 1972.6763008008008u,0 1973.6528408408408u,0 1973.653840840841u,1.5 1974.630380880881u,1.5 1974.6313808808811u,0 1975.6079209209206u,0 1975.6089209209208u,1.5 1976.5854609609607u,1.5 1976.586460960961u,0 1978.540541041041u,0 1978.5415410410412u,1.5 1979.5180810810812u,1.5 1979.5190810810814u,0 1982.4507012012011u,0 1982.4517012012013u,1.5 1983.4282412412413u,1.5 1983.4292412412415u,0 1988.3159414414415u,0 1988.3169414414417u,1.5 1989.2934814814816u,1.5 1989.2944814814819u,0 1995.1587217217213u,0 1995.1597217217216u,1.5 1996.1362617617615u,1.5 1996.1372617617617u,0 1997.1138018018016u,0 1997.1148018018018u,1.5 1999.068881881882u,1.5 1999.069881881882u,0 2002.979042042042u,0 2002.9800420420422u,1.5 2003.9565820820822u,1.5 2003.9575820820824u,0 2005.911662162162u,0 2005.9126621621622u,1.5 2006.8892022022021u,1.5 2006.8902022022023u,0 2017.6421426426425u,0 2017.6431426426427u,1.5 2018.6196826826827u,1.5 2018.6206826826829u,0 2020.5747627627625u,0 2020.5757627627627u,1.5 2021.5523028028026u,1.5 2021.5533028028028u,0 2024.4849229229226u,0 2024.4859229229228u,1.5 2025.4624629629627u,1.5 2025.463462962963u,0 2027.417543043043u,0 2027.4185430430432u,1.5 2030.350163163163u,1.5 2030.3511631631632u,0 2031.327703203203u,0 2031.3287032032033u,1.5 2032.3052432432432u,1.5 2032.3062432432434u,0 2033.2827832832834u,0 2033.2837832832836u,1.5 2038.1704834834836u,1.5 2038.1714834834838u,0 2039.1480235235233u,0 2039.1490235235235u,1.5 2045.9908038038036u,1.5 2045.9918038038038u,0 2046.9683438438437u,0 2046.969343843844u,1.5 2049.900963963964u,1.5 2049.901963963964u,0 2050.878504004004u,0 2050.879504004004u,1.5 2053.811124124124u,1.5 2053.8121241241242u,0 2058.698824324324u,0 2058.6998243243243u,1.5 2059.676364364364u,1.5 2059.677364364364u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2065.5416046046043u,1.5 2065.5426046046045u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2069.4517647647644u,0 2069.4527647647647u,1.5 2072.384384884885u,1.5 2072.3853848848853u,0 2074.339464964965u,0 2074.340464964965u,1.5 2076.294545045045u,1.5 2076.2955450450454u,0 2077.272085085085u,0 2077.2730850850853u,1.5 2078.249625125125u,1.5 2078.250625125125u,0 2088.025025525525u,0 2088.0260255255253u,1.5 2095.8453458458457u,1.5 2095.846345845846u,0 2097.8004259259255u,0 2097.8014259259257u,1.5 2098.777965965966u,1.5 2098.778965965966u,0 2099.755506006006u,0 2099.756506006006u,1.5 2100.733046046046u,1.5 2100.7340460460464u,0 2103.665666166166u,0 2103.666666166166u,1.5 2107.575826326326u,1.5 2107.576826326326u,0 2108.553366366366u,0 2108.554366366366u,1.5 2111.4859864864866u,1.5 2111.486986486487u,0 2115.3961466466467u,0 2115.397146646647u,1.5 2117.3512267267265u,1.5 2117.3522267267267u,0 2122.2389269269265u,0 2122.2399269269267u,1.5 2123.216466966967u,1.5 2123.217466966967u,0 2127.126627127127u,0 2127.127627127127u,1.5 2128.104167167167u,1.5 2128.105167167167u,0 2129.081707207207u,0 2129.082707207207u,1.5 2130.059247247247u,1.5 2130.0602472472474u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2138.8571076076073u,1.5 2138.8581076076075u,0 2139.8346476476477u,0 2139.835647647648u,1.5 2142.7672677677674u,1.5 2142.7682677677676u,0 2143.744807807808u,0 2143.745807807808u,1.5 2144.7223478478477u,1.5 2144.723347847848u,0 2147.654967967968u,0 2147.655967967968u,1.5 2148.632508008008u,1.5 2148.633508008008u,0 2149.610048048048u,0 2149.6110480480484u,1.5 2156.4528283283285u,1.5 2156.4538283283287u,0 2157.430368368368u,0 2157.431368368368u,1.5 2158.4079084084083u,1.5 2158.4089084084085u,0 2159.385448448448u,0 2159.3864484484484u,1.5 2160.3629884884886u,1.5 2160.3639884884888u,0 2161.3405285285285u,0 2161.3415285285287u,1.5 2166.228228728729u,1.5 2166.229228728729u,0 2168.1833088088088u,0 2168.184308808809u,1.5 2169.1608488488487u,1.5 2169.161848848849u,0 2171.115928928929u,0 2171.116928928929u,1.5 2173.071009009009u,1.5 2173.072009009009u,0 2175.026089089089u,0 2175.0270890890893u,1.5 2177.9587092092092u,1.5 2177.9597092092094u,0 2178.936249249249u,0 2178.9372492492494u,1.5 2179.913789289289u,1.5 2179.9147892892893u,0 2180.8913293293294u,0 2180.8923293293296u,1.5 2181.868869369369u,1.5 2181.869869369369u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2189.6891896896896u,1.5 2189.6901896896898u,0 2190.66672972973u,0 2190.66772972973u,1.5 2191.6442697697694u,1.5 2191.6452697697696u,0 2196.53196996997u,0 2196.53296996997u,1.5 2198.48705005005u,1.5 2198.4880500500503u,0 2199.46459009009u,0 2199.4655900900902u,1.5 2200.4421301301304u,1.5 2200.4431301301306u,0 2203.37475025025u,0 2203.3757502502503u,1.5 2204.35229029029u,1.5 2204.3532902902903u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2211.1950705705704u,1.5 2211.1960705705706u,0 2212.1726106106103u,0 2212.1736106106105u,1.5 2213.1501506506506u,1.5 2213.151150650651u,0 2215.105230730731u,0 2215.106230730731u,1.5 2216.0827707707704u,1.5 2216.0837707707706u,0 2219.015390890891u,0 2219.016390890891u,1.5 2222.925551051051u,1.5 2222.9265510510513u,0 2223.903091091091u,0 2223.9040910910912u,1.5 2224.8806311311314u,1.5 2224.8816311311316u,0 2225.858171171171u,0 2225.859171171171u,1.5 2226.835711211211u,1.5 2226.8367112112114u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2232.700951451451u,1.5 2232.7019514514514u,0 2242.4763518518516u,0 2242.477351851852u,1.5 2244.431431931932u,1.5 2244.432431931932u,0 2245.408971971972u,0 2245.409971971972u,1.5 2246.3865120120117u,1.5 2246.387512012012u,0 2250.296672172172u,0 2250.297672172172u,1.5 2255.184372372372u,1.5 2255.185372372372u,0 2256.161912412412u,0 2256.1629124124124u,1.5 2257.139452452452u,1.5 2257.1404524524523u,0 2258.1169924924925u,0 2258.1179924924927u,1.5 2259.0945325325324u,1.5 2259.0955325325326u,0 2261.0496126126122u,0 2261.0506126126124u,1.5 2262.0271526526526u,1.5 2262.028152652653u,0 2263.0046926926925u,0 2263.0056926926927u,1.5 2263.982232732733u,1.5 2263.983232732733u,0 2264.9597727727723u,0 2264.9607727727725u,1.5 2265.9373128128127u,1.5 2265.938312812813u,0 2266.9148528528526u,0 2266.915852852853u,1.5 2267.892392892893u,1.5 2267.893392892893u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2271.802553053053u,1.5 2271.8035530530533u,0 2272.780093093093u,0 2272.781093093093u,1.5 2274.735173173173u,1.5 2274.736173173173u,0 2275.712713213213u,0 2275.7137132132134u,1.5 2276.690253253253u,1.5 2276.6912532532533u,0 2281.577953453453u,0 2281.5789534534533u,1.5 2285.488113613613u,1.5 2285.4891136136134u,0 2286.4656536536536u,0 2286.466653653654u,1.5 2287.4431936936935u,1.5 2287.4441936936937u,0 2288.420733733734u,0 2288.421733733734u,1.5 2289.3982737737733u,1.5 2289.3992737737735u,0 2291.3533538538536u,0 2291.354353853854u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2294.285973973974u,0 2294.286973973974u,1.5 2295.2635140140137u,1.5 2295.264514014014u,0 2296.241054054054u,0 2296.2420540540543u,1.5 2297.218594094094u,1.5 2297.219594094094u,0 2298.1961341341344u,0 2298.1971341341346u,1.5 2299.173674174174u,1.5 2299.174674174174u,0 2304.0613743743743u,0 2304.0623743743745u,1.5 2307.9715345345344u,1.5 2307.9725345345346u,0 2308.9490745745743u,0 2308.9500745745745u,1.5 2309.926614614614u,1.5 2309.9276146146144u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2317.746934934935u,1.5 2317.747934934935u,0 2319.7020150150147u,0 2319.703015015015u,1.5 2320.679555055055u,1.5 2320.6805550550553u,0 2326.5447952952954u,0 2326.5457952952956u,1.5 2329.477415415415u,1.5 2329.4784154154154u,0 2330.454955455455u,0 2330.4559554554553u,1.5 2331.4324954954955u,1.5 2331.4334954954957u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2343.1629759759758u,1.5 2343.163975975976u,0 2344.1405160160157u,0 2344.141516016016u,1.5 2346.095596096096u,1.5 2346.096596096096u,0 2347.0731361361363u,0 2347.0741361361365u,1.5 2349.028216216216u,1.5 2349.0292162162164u,0 2350.9832962962964u,0 2350.9842962962966u,1.5 2353.915916416416u,1.5 2353.9169164164164u,0 2355.8709964964964u,0 2355.8719964964966u,1.5 2356.8485365365364u,1.5 2356.8495365365366u,0 2357.8260765765763u,0 2357.8270765765765u,1.5 2359.7811566566565u,1.5 2359.7821566566568u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2361.736236736737u,1.5 2361.737236736737u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2365.646396896897u,0 2365.647396896897u,1.5 2368.5790170170167u,1.5 2368.580017017017u,0 2369.556557057057u,0 2369.5575570570572u,1.5 2370.534097097097u,1.5 2370.535097097097u,0 2371.5116371371373u,0 2371.5126371371375u,1.5 2372.4891771771768u,1.5 2372.490177177177u,0 2378.354417417417u,0 2378.3554174174174u,1.5 2379.331957457457u,1.5 2379.3329574574573u,0 2380.3094974974974u,0 2380.3104974974976u,1.5 2386.174737737738u,1.5 2386.175737737738u,0 2387.1522777777777u,0 2387.153277777778u,1.5 2390.084897897898u,1.5 2390.085897897898u,0 2392.039977977978u,0 2392.0409779779784u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2394.972598098098u,0 2394.973598098098u,1.5 2395.9501381381383u,1.5 2395.9511381381385u,0 2397.905218218218u,0 2397.9062182182183u,1.5 2398.882758258258u,1.5 2398.8837582582582u,0 2400.8378383383383u,0 2400.8388383383385u,1.5 2402.792918418418u,1.5 2402.7939184184183u,0 2403.7704584584585u,0 2403.7714584584587u,1.5 2404.7479984984984u,1.5 2404.7489984984986u,0 2406.7030785785787u,0 2406.704078578579u,1.5 2407.680618618618u,1.5 2407.6816186186184u,0 2408.6581586586585u,0 2408.6591586586587u,1.5 2409.6356986986984u,1.5 2409.6366986986986u,0 2413.5458588588585u,0 2413.5468588588587u,1.5 2419.411099099099u,1.5 2419.412099099099u,0 2420.3886391391393u,0 2420.3896391391395u,1.5 2423.321259259259u,1.5 2423.322259259259u,0 2426.2538793793797u,0 2426.25487937938u,1.5 2427.231419419419u,1.5 2427.2324194194193u,0 2430.1640395395393u,0 2430.1650395395395u,1.5 2432.119119619619u,1.5 2432.1201196196193u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.0068198198196u,1.5 2437.00781981982u,0 2438.9618998999u,0 2438.9628998999u,1.5 2446.78222022022u,1.5 2446.7832202202203u,0 2447.75976026026u,0 2447.76076026026u,1.5 2449.7148403403403u,1.5 2449.7158403403405u,0 2451.66992042042u,0 2451.6709204204203u,1.5 2452.6474604604605u,1.5 2452.6484604604607u,0 2453.6250005005004u,0 2453.6260005005006u,1.5 2454.6025405405403u,1.5 2454.6035405405405u,0 2463.400400900901u,0 2463.401400900901u,1.5 2465.355480980981u,1.5 2465.3564809809814u,0 2466.3330210210206u,0 2466.334021021021u,1.5 2467.310561061061u,1.5 2467.311561061061u,0 2469.2656411411413u,0 2469.2666411411415u,1.5 2470.243181181181u,1.5 2470.2441811811814u,0 2472.198261261261u,0 2472.199261261261u,1.5 2473.1758013013014u,1.5 2473.1768013013016u,0 2475.1308813813816u,0 2475.131881381382u,1.5 2476.108421421421u,1.5 2476.1094214214213u,0 2477.0859614614615u,0 2477.0869614614617u,1.5 2479.0410415415413u,1.5 2479.0420415415415u,0 2480.996121621621u,0 2480.9971216216213u,1.5 2484.9062817817817u,1.5 2484.907281781782u,0 2485.8838218218216u,0 2485.884821821822u,1.5 2487.838901901902u,1.5 2487.839901901902u,0 2489.793981981982u,0 2489.7949819819823u,1.5 2494.681682182182u,1.5 2494.6826821821824u,0 2495.659222222222u,0 2495.6602222222223u,1.5 2502.5020025025024u,1.5 2502.5030025025026u,0 2505.434622622622u,0 2505.4356226226223u,1.5 2507.3897027027024u,1.5 2507.3907027027026u,0 2508.3672427427427u,0 2508.368242742743u,1.5 2511.2998628628625u,1.5 2511.3008628628627u,0 2512.277402902903u,0 2512.278402902903u,1.5 2513.2549429429428u,1.5 2513.255942942943u,0 2516.187563063063u,0 2516.188563063063u,1.5 2522.0528033033033u,1.5 2522.0538033033035u,0 2523.0303433433432u,0 2523.0313433433435u,1.5 2524.0078833833836u,1.5 2524.008883383384u,0 2524.985423423423u,0 2524.9864234234233u,1.5 2526.9405035035034u,1.5 2526.9415035035036u,0 2527.9180435435437u,0 2527.919043543544u,1.5 2528.8955835835836u,1.5 2528.896583583584u,0 2530.8506636636635u,0 2530.8516636636637u,1.5 2531.8282037037034u,1.5 2531.8292037037036u,0 2532.8057437437437u,0 2532.806743743744u,1.5 2533.7832837837836u,1.5 2533.784283783784u,0 2535.7383638638635u,0 2535.7393638638637u,1.5 2536.715903903904u,1.5 2536.716903903904u,0 2538.670983983984u,0 2538.6719839839843u,1.5 2539.6485240240236u,1.5 2539.649524024024u,0 2540.626064064064u,0 2540.627064064064u,1.5 2542.581144144144u,1.5 2542.5821441441444u,0 2545.513764264264u,0 2545.514764264264u,1.5 2546.4913043043043u,1.5 2546.4923043043045u,0 2549.423924424424u,0 2549.4249244244243u,1.5 2550.4014644644644u,1.5 2550.4024644644646u,0 2552.3565445445447u,0 2552.357544544545u,1.5 2556.2667047047044u,1.5 2556.2677047047046u,0 2557.2442447447447u,0 2557.245244744745u,1.5 2559.1993248248245u,1.5 2559.2003248248247u,0 2560.1768648648645u,0 2560.1778648648647u,1.5 2563.109484984985u,1.5 2563.1104849849853u,0 2564.0870250250246u,0 2564.0880250250248u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2572.8848853853856u,1.5 2572.885885385386u,0 2574.8399654654654u,0 2574.8409654654656u,1.5 2575.8175055055053u,1.5 2575.8185055055055u,0 2577.7725855855856u,0 2577.773585585586u,1.5 2579.7276656656654u,1.5 2579.7286656656656u,0 2582.6602857857856u,0 2582.661285785786u,1.5 2583.6378258258255u,1.5 2583.6388258258257u,0 2584.6153658658654u,0 2584.6163658658656u,1.5 2588.5255260260255u,1.5 2588.5265260260257u,0 2590.480606106106u,0 2590.481606106106u,1.5 2593.413226226226u,1.5 2593.414226226226u,0 2594.390766266266u,0 2594.391766266266u,1.5 2595.3683063063063u,1.5 2595.3693063063065u,0 2597.3233863863866u,0 2597.324386386387u,1.5 2598.300926426426u,1.5 2598.3019264264262u,0 2599.2784664664664u,0 2599.2794664664666u,1.5 2600.2560065065063u,1.5 2600.2570065065065u,0 2602.2110865865866u,0 2602.212086586587u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2607.0987867867866u,1.5 2607.099786786787u,0 2613.941567067067u,0 2613.942567067067u,1.5 2617.851727227227u,1.5 2617.852727227227u,0 2618.829267267267u,0 2618.830267267267u,1.5 2620.784347347347u,1.5 2620.7853473473474u,0 2623.7169674674674u,0 2623.7179674674676u,1.5 2627.6271276276275u,1.5 2627.6281276276277u,0 2630.5597477477477u,0 2630.560747747748u,1.5 2636.424987987988u,1.5 2636.4259879879883u,0 2638.380068068068u,0 2638.381068068068u,1.5 2639.357608108108u,1.5 2639.358608108108u,0 2643.267768268268u,0 2643.268768268268u,1.5 2648.1554684684684u,1.5 2648.1564684684686u,0 2649.1330085085083u,0 2649.1340085085085u,1.5 2650.1105485485486u,1.5 2650.111548548549u,0 2652.065628628629u,0 2652.066628628629u,1.5 2653.0431686686684u,1.5 2653.0441686686686u,0 2654.0207087087088u,0 2654.021708708709u,1.5 2654.9982487487487u,1.5 2654.999248748749u,0 2655.9757887887886u,0 2655.976788788789u,1.5 2656.953328828829u,1.5 2656.954328828829u,0 2657.9308688688684u,0 2657.9318688688686u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2668.6838093093093u,0 2668.6848093093095u,1.5 2673.5715095095093u,1.5 2673.5725095095095u,0 2674.5490495495496u,0 2674.55004954955u,1.5 2676.50412962963u,1.5 2676.50512962963u,0 2677.4816696696694u,0 2677.4826696696696u,1.5 2678.4592097097097u,1.5 2678.46020970971u,0 2679.4367497497497u,0 2679.43774974975u,1.5 2680.4142897897896u,1.5 2680.4152897897898u,0 2681.39182982983u,0 2681.39282982983u,1.5 2686.27953003003u,1.5 2686.28053003003u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2689.21215015015u,0 2689.2131501501503u,1.5 2690.18969019019u,1.5 2690.1906901901903u,0 2692.14477027027u,0 2692.14577027027u,1.5 2694.09985035035u,1.5 2694.1008503503504u,0 2695.0773903903905u,0 2695.0783903903907u,1.5 2698.0100105105103u,1.5 2698.0110105105105u,0 2698.9875505505506u,0 2698.988550550551u,1.5 2699.9650905905905u,1.5 2699.9660905905907u,0 2700.942630630631u,0 2700.943630630631u,1.5 2701.9201706706704u,1.5 2701.9211706706706u,0 2702.8977107107107u,0 2702.898710710711u,1.5 2704.8527907907906u,1.5 2704.8537907907908u,0 2705.830330830831u,0 2705.831330830831u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2708.7629509509507u,0 2708.763950950951u,1.5 2709.740490990991u,1.5 2709.741490990991u,0 2710.718031031031u,0 2710.719031031031u,1.5 2711.695571071071u,1.5 2711.696571071071u,0 2712.6731111111108u,0 2712.674111111111u,1.5 2713.650651151151u,1.5 2713.6516511511513u,0 2714.628191191191u,0 2714.6291911911912u,1.5 2716.583271271271u,1.5 2716.584271271271u,0 2718.538351351351u,0 2718.5393513513513u,1.5 2719.5158913913915u,1.5 2719.5168913913917u,0 2721.4709714714713u,0 2721.4719714714715u,1.5 2723.4260515515516u,1.5 2723.427051551552u,0 2724.4035915915915u,0 2724.4045915915917u,1.5 2725.381131631632u,1.5 2725.382131631632u,0 2727.3362117117117u,0 2727.337211711712u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2732.2239119119117u,1.5 2732.224911911912u,0 2737.1116121121117u,0 2737.112612112112u,1.5 2739.066692192192u,1.5 2739.067692192192u,0 2740.0442322322324u,0 2740.0452322322326u,1.5 2741.021772272272u,1.5 2741.022772272272u,0 2745.9094724724723u,0 2745.9104724724725u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2755.6848728728723u,0 2755.6858728728726u,1.5 2757.6399529529526u,1.5 2757.640952952953u,0 2759.595033033033u,0 2759.596033033033u,1.5 2760.572573073073u,1.5 2760.573573073073u,0 2763.505193193193u,0 2763.506193193193u,1.5 2765.460273273273u,1.5 2765.461273273273u,0 2766.437813313313u,0 2766.4388133133134u,1.5 2768.3928933933935u,1.5 2768.3938933933937u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2775.2356736736733u,0 2775.2366736736735u,1.5 2777.1907537537536u,1.5 2777.191753753754u,0 2778.168293793794u,0 2778.169293793794u,1.5 2782.0784539539536u,1.5 2782.079453953954u,0 2785.9886141141137u,0 2785.989614114114u,1.5 2786.966154154154u,1.5 2786.9671541541543u,0 2787.943694194194u,0 2787.944694194194u,1.5 2790.876314314314u,1.5 2790.8773143143144u,0 2791.853854354354u,0 2791.8548543543543u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2793.8089344344344u,0 2793.8099344344346u,1.5 2794.7864744744743u,1.5 2794.7874744744745u,0 2795.764014514514u,0 2795.7650145145144u,1.5 2796.7415545545546u,1.5 2796.7425545545548u,0 2797.7190945945945u,0 2797.7200945945947u,1.5 2804.561874874875u,1.5 2804.562874874875u,0 2807.494494994995u,0 2807.495494994995u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2822.1575955955955u,0 2822.1585955955957u,1.5 2828.022835835836u,1.5 2828.023835835836u,0 2830.9554559559556u,0 2830.956455955956u,1.5 2831.932995995996u,1.5 2831.933995995996u,0 2832.910536036036u,0 2832.911536036036u,1.5 2833.888076076076u,1.5 2833.889076076076u,0 2834.8656161161157u,0 2834.866616116116u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2841.7083963963964u,0 2841.7093963963966u,1.5 2842.6859364364364u,1.5 2842.6869364364366u,0 2844.641016516516u,0 2844.6420165165164u,1.5 2845.6185565565565u,1.5 2845.6195565565567u,0 2849.5287167167166u,0 2849.529716716717u,1.5 2850.5062567567566u,1.5 2850.5072567567568u,0 2851.483796796797u,0 2851.484796796797u,1.5 2852.461336836837u,1.5 2852.462336836837u,0 2856.371496996997u,0 2856.372496996997u,1.5 2857.349037037037u,1.5 2857.350037037037u,0 2858.3265770770768u,0 2858.327577077077u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2864.191817317317u,1.5 2864.1928173173173u,0 2868.1019774774772u,0 2868.1029774774775u,1.5 2869.079517517517u,1.5 2869.0805175175174u,0 2870.0570575575575u,0 2870.0580575575577u,1.5 2871.0345975975974u,1.5 2871.0355975975976u,0 2872.012137637638u,0 2872.013137637638u,1.5 2876.899837837838u,1.5 2876.900837837838u,0 2877.877377877878u,0 2877.8783778778784u,1.5 2878.8549179179176u,1.5 2878.855917917918u,0 2880.809997997998u,0 2880.810997997998u,1.5 2883.7426181181177u,1.5 2883.743618118118u,0 2885.697698198198u,0 2885.698698198198u,1.5 2886.6752382382383u,1.5 2886.6762382382385u,0 2887.652778278278u,0 2887.6537782782784u,1.5 2888.630318318318u,1.5 2888.6313183183183u,0 2891.5629384384383u,0 2891.5639384384385u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2897.4281786786787u,0 2897.429178678679u,1.5 2898.4057187187186u,1.5 2898.406718718719u,0 2901.338338838839u,0 2901.339338838839u,1.5 2906.226039039039u,1.5 2906.227039039039u,0 2908.1811191191186u,0 2908.182119119119u,1.5 2911.1137392392393u,1.5 2911.1147392392395u,0 2912.091279279279u,0 2912.0922792792794u,1.5 2913.068819319319u,1.5 2913.0698193193193u,0 2917.956519519519u,0 2917.9575195195193u,1.5 2920.88913963964u,1.5 2920.89013963964u,0 2921.8666796796797u,0 2921.86767967968u,1.5 2922.8442197197196u,1.5 2922.84521971972u,0 2923.8217597597595u,0 2923.8227597597597u,1.5 2925.77683983984u,1.5 2925.77783983984u,0 2926.75437987988u,0 2926.7553798798804u,1.5 2927.7319199199196u,1.5 2927.73291991992u,0 2929.687u,0 2929.688u,1.5 2931.64208008008u,1.5 2931.6430800800804u,0 2932.6196201201196u,0 2932.62062012012u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2936.52978028028u,0 2936.5307802802804u,1.5 2937.50732032032u,1.5 2937.5083203203203u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2942.39502052052u,0 2942.3960205205203u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 2948.2602607607605u,0 2948.2612607607607u,1.5 2949.237800800801u,1.5 2949.238800800801u,0 2950.215340840841u,0 2950.216340840841u,1.5 2952.1704209209206u,1.5 2952.171420920921u,0 2953.147960960961u,0 2953.148960960961u,1.5 2955.103041041041u,1.5 2955.104041041041u,0 2957.0581211211206u,0 2957.059121121121u,1.5 2958.035661161161u,1.5 2958.036661161161u,0 2959.013201201201u,0 2959.014201201201u,1.5 2960.968281281281u,1.5 2960.9692812812814u,0 2966.833521521521u,0 2966.8345215215213u,1.5 2967.8110615615615u,1.5 2967.8120615615617u,0 2968.7886016016014u,0 2968.7896016016016u,1.5 2969.7661416416418u,1.5 2969.767141641642u,0 2970.7436816816817u,0 2970.744681681682u,1.5 2972.6987617617615u,1.5 2972.6997617617617u,0 2974.6538418418418u,0 2974.654841841842u,1.5 2975.631381881882u,1.5 2975.6323818818823u,0 2980.519082082082u,0 2980.5200820820824u,1.5 2981.4966221221216u,1.5 2981.497622122122u,0 2983.451702202202u,0 2983.452702202202u,1.5 2984.4292422422423u,1.5 2984.4302422422425u,0 2986.384322322322u,0 2986.3853223223223u,1.5 2988.3394024024024u,1.5 2988.3404024024026u,0 2989.3169424424423u,0 2989.3179424424425u,1.5 2990.2944824824826u,1.5 2990.295482482483u,0 2993.2271026026024u,0 2993.2281026026026u,1.5 2994.2046426426427u,1.5 2994.205642642643u,0 2997.1372627627625u,0 2997.1382627627627u,1.5 2998.114802802803u,1.5 2998.115802802803u,0 2999.0923428428428u,0 2999.093342842843u,1.5 3000.069882882883u,1.5 3000.0708828828833u,0 3003.980043043043u,0 3003.9810430430434u,1.5 3004.957583083083u,1.5 3004.9585830830833u,0 3010.822823323323u,0 3010.8238233233233u,1.5 3011.800363363363u,1.5 3011.801363363363u,0 3014.7329834834836u,0 3014.733983483484u,1.5 3015.710523523523u,1.5 3015.7115235235233u,0 3017.6656036036034u,0 3017.6666036036036u,1.5 3018.6431436436437u,1.5 3018.644143643644u,0 3022.553303803804u,0 3022.554303803804u,1.5 3023.5308438438437u,1.5 3023.531843843844u,0 3026.463463963964u,0 3026.464463963964u,1.5 3027.441004004004u,1.5 3027.442004004004u,0 3028.418544044044u,0 3028.4195440440444u,1.5 3029.396084084084u,1.5 3029.3970840840843u,0 3030.373624124124u,0 3030.3746241241242u,1.5 3032.328704204204u,1.5 3032.329704204204u,0 3033.306244244244u,0 3033.3072442442444u,1.5 3036.238864364364u,1.5 3036.239864364364u,0 3037.2164044044043u,0 3037.2174044044045u,1.5 3039.1714844844846u,1.5 3039.172484484485u,0 3040.149024524524u,0 3040.1500245245243u,1.5 3043.0816446446447u,1.5 3043.082644644645u,0 3044.0591846846846u,0 3044.060184684685u,1.5 3046.0142647647644u,1.5 3046.0152647647647u,0 3046.991804804805u,0 3046.992804804805u,1.5 3048.946884884885u,1.5 3048.9478848848853u,0 3050.901964964965u,0 3050.902964964965u,1.5 3051.879505005005u,1.5 3051.880505005005u,0 3059.699825325325u,0 3059.7008253253252u,1.5 3061.6549054054053u,1.5 3061.6559054054055u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3064.587525525525u,1.5 3064.5885255255253u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3069.4752257257255u,1.5 3069.4762257257257u,0 3070.4527657657654u,0 3070.4537657657656u,1.5 3073.385385885886u,1.5 3073.3863858858863u,0 3076.318006006006u,0 3076.319006006006u,1.5 3077.295546046046u,1.5 3077.2965460460464u,0 3081.205706206206u,0 3081.206706206206u,1.5 3082.183246246246u,1.5 3082.1842462462464u,0 3085.115866366366u,0 3085.116866366366u,1.5 3086.0934064064063u,1.5 3086.0944064064065u,0 3089.026026526526u,0 3089.0270265265262u,1.5 3093.9137267267265u,1.5 3093.9147267267267u,0 3094.8912667667664u,0 3094.8922667667666u,1.5 3096.8463468468467u,1.5 3096.847346846847u,0 3097.823886886887u,0 3097.8248868868873u,1.5 3100.756507007007u,1.5 3100.757507007007u,0 3102.711587087087u,0 3102.7125870870873u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3108.576827327327u,1.5 3108.577827327327u,0 3109.554367367367u,0 3109.555367367367u,1.5 3112.4869874874876u,1.5 3112.4879874874878u,0 3113.464527527527u,0 3113.4655275275272u,1.5 3114.4420675675674u,1.5 3114.4430675675676u,0 3119.3297677677674u,0 3119.3307677677676u,1.5 3121.2848478478477u,1.5 3121.285847847848u,0 3122.262387887888u,0 3122.2633878878883u,1.5 3128.127628128128u,1.5 3128.128628128128u,0 3129.105168168168u,0 3129.106168168168u,1.5 3130.0827082082083u,1.5 3130.0837082082085u,0 3132.037788288288u,0 3132.0387882882883u,1.5 3133.992868368368u,1.5 3133.993868368368u,0 3134.9704084084083u,0 3134.9714084084085u,1.5 3136.9254884884886u,1.5 3136.9264884884888u,0 3137.9030285285285u,0 3137.9040285285287u,1.5 3139.8581086086083u,1.5 3139.8591086086085u,0 3140.8356486486487u,0 3140.836648648649u,1.5 3141.8131886886886u,1.5 3141.814188688689u,0 3142.790728728729u,0 3142.791728728729u,1.5 3143.7682687687684u,1.5 3143.7692687687686u,0 3144.7458088088088u,0 3144.746808808809u,1.5 3146.700888888889u,1.5 3146.7018888888892u,0 3147.678428928929u,0 3147.679428928929u,1.5 3148.655968968969u,1.5 3148.656968968969u,0 3149.633509009009u,0 3149.634509009009u,1.5 3151.588589089089u,1.5 3151.5895890890893u,0 3153.543669169169u,0 3153.544669169169u,1.5 3154.5212092092092u,1.5 3154.5222092092094u,0 3155.498749249249u,0 3155.4997492492494u,1.5 3157.4538293293294u,1.5 3157.4548293293296u,0 3160.386449449449u,0 3160.3874494494494u,1.5 3162.3415295295295u,1.5 3162.3425295295297u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3164.2966096096093u,1.5 3164.2976096096095u,0 3166.2516896896896u,0 3166.2526896896898u,1.5 3168.2067697697694u,1.5 3168.2077697697696u,0 3169.1843098098097u,0 3169.18530980981u,1.5 3170.1618498498497u,1.5 3170.16284984985u,0 3174.0720100100098u,0 3174.07301001001u,1.5 3175.04955005005u,1.5 3175.0505500500503u,0 3176.02709009009u,0 3176.0280900900902u,1.5 3177.98217017017u,1.5 3177.98317017017u,0 3178.9597102102102u,0 3178.9607102102104u,1.5 3179.93725025025u,1.5 3179.9382502502503u,0 3180.91479029029u,0 3180.9157902902903u,1.5 3181.8923303303304u,1.5 3181.8933303303306u,0 3183.8474104104102u,0 3183.8484104104105u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3187.7575705705704u,0 3187.7585705705706u,1.5 3190.6901906906905u,1.5 3190.6911906906907u,0 3191.667730730731u,0 3191.668730730731u,1.5 3192.6452707707704u,1.5 3192.6462707707706u,0 3195.577890890891u,0 3195.578890890891u,1.5 3196.555430930931u,1.5 3196.556430930931u,0 3197.532970970971u,0 3197.533970970971u,1.5 3203.398211211211u,1.5 3203.3992112112114u,0 3204.375751251251u,0 3204.3767512512513u,1.5 3205.353291291291u,1.5 3205.3542912912912u,0 3209.263451451451u,0 3209.2644514514514u,1.5 3213.1736116116112u,1.5 3213.1746116116115u,0 3214.1511516516516u,0 3214.152151651652u,1.5 3217.0837717717714u,1.5 3217.0847717717716u,0 3218.0613118118117u,0 3218.062311811812u,1.5 3219.0388518518516u,1.5 3219.039851851852u,0 3220.016391891892u,0 3220.017391891892u,1.5 3223.926552052052u,1.5 3223.9275520520523u,0 3224.904092092092u,0 3224.905092092092u,1.5 3225.8816321321324u,1.5 3225.8826321321326u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3234.6794924924925u,1.5 3234.6804924924927u,0 3238.5896526526526u,0 3238.590652652653u,1.5 3240.544732732733u,1.5 3240.545732732733u,0 3241.5222727727723u,0 3241.5232727727725u,1.5 3244.454892892893u,1.5 3244.455892892893u,0 3246.409972972973u,0 3246.410972972973u,1.5 3247.3875130130127u,1.5 3247.388513013013u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3254.2302932932935u,1.5 3254.2312932932937u,0 3261.0730735735733u,0 3261.0740735735735u,1.5 3262.050613613613u,1.5 3262.0516136136134u,0 3263.0281536536536u,0 3263.029153653654u,1.5 3264.983233733734u,1.5 3264.984233733734u,0 3266.9383138138137u,0 3266.939313813814u,1.5 3267.9158538538536u,1.5 3267.916853853854u,0 3269.870933933934u,0 3269.871933933934u,1.5 3270.848473973974u,1.5 3270.849473973974u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3273.781094094094u,0 3273.782094094094u,1.5 3276.713714214214u,1.5 3276.7147142142144u,0 3280.6238743743743u,0 3280.6248743743745u,1.5 3281.601414414414u,1.5 3281.6024144144144u,0 3283.5564944944945u,0 3283.5574944944947u,1.5 3287.4666546546546u,1.5 3287.467654654655u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3297.242055055055u,1.5 3297.2430550550553u,0 3298.219595095095u,0 3298.220595095095u,1.5 3299.1971351351353u,1.5 3299.1981351351355u,0 3300.174675175175u,0 3300.175675175175u,1.5 3306.039915415415u,1.5 3306.0409154154154u,0 3307.017455455455u,0 3307.0184554554553u,1.5 3307.9949954954955u,1.5 3307.9959954954957u,0 3309.9500755755753u,0 3309.9510755755755u,1.5 3310.927615615615u,1.5 3310.9286156156154u,0 3312.8826956956955u,0 3312.8836956956957u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3315.8153158158157u,0 3315.816315815816u,1.5 3317.770395895896u,1.5 3317.771395895896u,0 3318.747935935936u,0 3318.748935935936u,1.5 3319.7254759759758u,1.5 3319.726475975976u,0 3323.6356361361363u,0 3323.6366361361365u,1.5 3324.613176176176u,1.5 3324.614176176176u,0 3325.590716216216u,0 3325.5917162162164u,1.5 3326.568256256256u,1.5 3326.5692562562563u,0 3330.478416416416u,0 3330.4794164164164u,1.5 3331.455956456456u,1.5 3331.4569564564563u,0 3332.4334964964964u,0 3332.4344964964966u,1.5 3333.4110365365364u,1.5 3333.4120365365366u,0 3335.366116616616u,0 3335.3671166166164u,1.5 3337.3211966966965u,1.5 3337.3221966966967u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3342.208896896897u,1.5 3342.209896896897u,0 3343.186436936937u,0 3343.187436936937u,1.5 3346.119057057057u,1.5 3346.1200570570572u,0 3350.029217217217u,0 3350.0302172172173u,1.5 3351.006757257257u,1.5 3351.0077572572573u,0 3351.9842972972974u,0 3351.9852972972976u,1.5 3355.894457457457u,1.5 3355.8954574574573u,0 3356.8719974974974u,0 3356.8729974974976u,1.5 3357.8495375375373u,1.5 3357.8505375375375u,0 3360.7821576576575u,0 3360.7831576576577u,1.5 3363.7147777777773u,1.5 3363.7157777777775u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3369.5800180180177u,1.5 3369.581018018018u,0 3371.535098098098u,0 3371.536098098098u,1.5 3372.5126381381383u,1.5 3372.5136381381385u,0 3373.4901781781778u,0 3373.491178178178u,1.5 3374.467718218218u,1.5 3374.4687182182183u,0 3379.355418418418u,0 3379.3564184184183u,1.5 3382.2880385385383u,1.5 3382.2890385385385u,0 3383.2655785785787u,0 3383.266578578579u,1.5 3386.1981986986984u,1.5 3386.1991986986986u,0 3387.175738738739u,0 3387.176738738739u,1.5 3390.1083588588585u,1.5 3390.1093588588587u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.0185190190186u,1.5 3394.019519019019u,0 3394.996059059059u,0 3394.997059059059u,1.5 3398.906219219219u,1.5 3398.9072192192193u,0 3399.883759259259u,0 3399.884759259259u,1.5 3400.8612992992994u,1.5 3400.8622992992996u,0 3401.8388393393393u,0 3401.8398393393395u,1.5 3403.793919419419u,1.5 3403.7949194194193u,0 3407.7040795795797u,0 3407.70507957958u,1.5 3409.6591596596595u,1.5 3409.6601596596597u,0 3410.6366996996994u,0 3410.6376996996996u,1.5 3411.61423973974u,1.5 3411.61523973974u,0 3412.5917797797797u,0 3412.59277977978u,1.5 3414.5468598598595u,1.5 3414.5478598598597u,0 3415.5243998999u,0 3415.5253998999u,1.5 3420.4121001001u,1.5 3420.4131001001u,0 3421.3896401401403u,0 3421.3906401401405u,1.5 3422.36718018018u,1.5 3422.3681801801804u,0 3424.32226026026u,0 3424.32326026026u,1.5 3425.2998003003004u,1.5 3425.3008003003006u,0 3427.2548803803807u,0 3427.255880380381u,1.5 3428.23242042042u,1.5 3428.2334204204203u,0 3429.2099604604605u,0 3429.2109604604607u,1.5 3430.1875005005004u,1.5 3430.1885005005006u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3437.0302807807807u,0 3437.031280780781u,1.5 3438.0078208208206u,1.5 3438.008820820821u,0 3438.9853608608605u,0 3438.9863608608607u,1.5 3446.805681181181u,1.5 3446.8066811811814u,0 3447.783221221221u,0 3447.7842212212213u,1.5 3450.7158413413413u,1.5 3450.7168413413415u,0 3452.670921421421u,0 3452.6719214214213u,1.5 3453.6484614614615u,1.5 3453.6494614614617u,0 3454.6260015015014u,0 3454.6270015015016u,1.5 3456.5810815815817u,1.5 3456.582081581582u,0 3460.4912417417418u,0 3460.492241741742u,1.5 3461.4687817817817u,1.5 3461.469781781782u,0 3465.378941941942u,0 3465.379941941942u,1.5 3466.356481981982u,1.5 3466.3574819819823u,0 3467.3340220220216u,0 3467.335022022022u,1.5 3468.311562062062u,1.5 3468.312562062062u,0 3469.289102102102u,0 3469.290102102102u,1.5 3470.2666421421422u,1.5 3470.2676421421424u,0 3472.221722222222u,0 3472.2227222222223u,1.5 3473.199262262262u,1.5 3473.200262262262u,0 3474.1768023023023u,0 3474.1778023023026u,1.5 3475.1543423423423u,1.5 3475.1553423423425u,0 3476.1318823823826u,0 3476.132882382383u,1.5 3478.0869624624625u,1.5 3478.0879624624627u,0 3479.0645025025024u,0 3479.0655025025026u,1.5 3481.0195825825826u,1.5 3481.020582582583u,0 3481.997122622622u,0 3481.9981226226223u,1.5 3482.9746626626625u,1.5 3482.9756626626627u,0 3483.9522027027024u,0 3483.9532027027026u,1.5 3493.727603103103u,1.5 3493.728603103103u,0 3494.7051431431432u,0 3494.7061431431434u,1.5 3495.682683183183u,1.5 3495.6836831831833u,0 3496.660223223223u,0 3496.6612232232233u,1.5 3501.547923423423u,1.5 3501.5489234234233u,0 3503.5030035035034u,0 3503.5040035035036u,1.5 3521.098724224224u,1.5 3521.0997242242242u,0 3522.076264264264u,0 3522.077264264264u,1.5 3525.0088843843846u,1.5 3525.009884384385u,0 3526.9639644644644u,0 3526.9649644644646u,1.5 3527.9415045045043u,1.5 3527.9425045045045u,0 3529.8965845845846u,0 3529.897584584585u,1.5 3530.8741246246245u,1.5 3530.8751246246247u,0 3531.8516646646644u,0 3531.8526646646646u,1.5 3533.8067447447447u,1.5 3533.807744744745u,0 3535.7618248248245u,0 3535.7628248248247u,1.5 3536.7393648648645u,1.5 3536.7403648648647u,0 3537.716904904905u,0 3537.717904904905u,1.5 3539.671984984985u,1.5 3539.6729849849853u,0 3540.6495250250246u,0 3540.6505250250248u,1.5 3541.627065065065u,1.5 3541.628065065065u,0 3542.604605105105u,0 3542.605605105105u,1.5 3543.582145145145u,1.5 3543.5831451451454u,0 3546.514765265265u,0 3546.515765265265u,1.5 3547.4923053053053u,1.5 3547.4933053053055u,0 3548.469845345345u,0 3548.4708453453454u,1.5 3549.4473853853856u,1.5 3549.448385385386u,0 3551.4024654654654u,0 3551.4034654654656u,1.5 3553.3575455455457u,1.5 3553.358545545546u,0 3554.3350855855856u,0 3554.336085585586u,1.5 3555.3126256256255u,1.5 3555.3136256256257u,0 3556.2901656656654u,0 3556.2911656656656u,1.5 3561.1778658658654u,1.5 3561.1788658658656u,0 3562.155405905906u,0 3562.156405905906u,1.5 3564.110485985986u,1.5 3564.1114859859863u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.998186186186u,0 3568.9991861861863u,1.5 3570.953266266266u,1.5 3570.954266266266u,0 3574.863426426426u,0 3574.8644264264262u,1.5 3576.8185065065063u,1.5 3576.8195065065065u,0 3577.7960465465467u,0 3577.797046546547u,1.5 3578.7735865865866u,1.5 3578.774586586587u,0 3579.7511266266265u,0 3579.7521266266267u,1.5 3581.7062067067063u,1.5 3581.7072067067065u,0 3582.6837467467467u,0 3582.684746746747u,1.5 3583.6612867867866u,1.5 3583.662286786787u,0 3584.6388268268265u,0 3584.6398268268267u,1.5 3586.593906906907u,1.5 3586.594906906907u,0 3588.548986986987u,0 3588.5499869869873u,1.5 3589.5265270270265u,1.5 3589.5275270270267u,0 3597.346847347347u,0 3597.3478473473474u,1.5 3598.3243873873876u,1.5 3598.3253873873878u,0 3599.301927427427u,0 3599.302927427427u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3609.0773278278275u,1.5 3609.0783278278277u,0 3612.0099479479477u,0 3612.010947947948u,1.5 3612.987487987988u,1.5 3612.9884879879883u,0 3613.9650280280275u,0 3613.9660280280277u,1.5 3615.920108108108u,1.5 3615.921108108108u,0 3616.897648148148u,0 3616.8986481481484u,1.5 3617.875188188188u,1.5 3617.8761881881883u,0 3619.830268268268u,0 3619.831268268268u,1.5 3621.785348348348u,1.5 3621.7863483483484u,0 3622.7628883883885u,0 3622.7638883883888u,1.5 3623.740428428428u,1.5 3623.741428428428u,0 3624.7179684684684u,0 3624.7189684684686u,1.5 3625.6955085085083u,1.5 3625.6965085085085u,0 3627.6505885885886u,0 3627.6515885885888u,1.5 3628.6281286286285u,1.5 3628.6291286286287u,0 3630.5832087087088u,0 3630.584208708709u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3640.358609109109u,0 3640.359609109109u,1.5 3641.336149149149u,1.5 3641.3371491491494u,0 3643.2912292292294u,0 3643.2922292292296u,1.5 3650.1340095095093u,1.5 3650.1350095095095u,0 3651.1115495495496u,0 3651.11254954955u,1.5 3652.0890895895895u,1.5 3652.0900895895898u,0 3655.9992497497497u,0 3656.00024974975u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3666.75219019019u,0 3666.7531901901903u,1.5 3667.7297302302304u,1.5 3667.7307302302306u,0 3670.66235035035u,0 3670.6633503503504u,1.5 3675.5500505505506u,1.5 3675.551050550551u,0 3676.5275905905905u,0 3676.5285905905907u,1.5 3677.505130630631u,1.5 3677.506130630631u,0 3678.4826706706704u,0 3678.4836706706706u,1.5 3679.4602107107107u,1.5 3679.461210710711u,0 3682.392830830831u,0 3682.393830830831u,1.5 3685.3254509509507u,1.5 3685.326450950951u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3689.2356111111108u,0 3689.236611111111u,1.5 3690.213151151151u,1.5 3690.2141511511513u,0 3691.190691191191u,0 3691.1916911911912u,1.5 3693.145771271271u,1.5 3693.146771271271u,0 3694.123311311311u,0 3694.1243113113114u,1.5 3697.0559314314314u,1.5 3697.0569314314316u,0 3698.0334714714713u,0 3698.0344714714715u,1.5 3699.0110115115112u,1.5 3699.0120115115114u,0 3702.9211716716713u,0 3702.9221716716715u,1.5 3703.8987117117117u,1.5 3703.899711711712u,0 3705.8537917917915u,0 3705.8547917917917u,1.5 3707.8088718718714u,1.5 3707.8098718718716u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3713.6741121121117u,0 3713.675112112112u,1.5 3718.561812312312u,1.5 3718.5628123123124u,0 3719.539352352352u,0 3719.5403523523523u,1.5 3720.5168923923925u,1.5 3720.5178923923927u,0 3723.4495125125122u,0 3723.4505125125124u,1.5 3725.4045925925925u,1.5 3725.4055925925927u,0 3726.382132632633u,0 3726.383132632633u,1.5 3728.3372127127127u,1.5 3728.338212712713u,0 3729.3147527527526u,0 3729.315752752753u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3732.2473728728723u,0 3732.2483728728726u,1.5 3735.179992992993u,1.5 3735.180992992993u,0 3736.157533033033u,0 3736.158533033033u,1.5 3740.067693193193u,1.5 3740.068693193193u,0 3744.9553933933935u,0 3744.9563933933937u,1.5 3745.9329334334334u,1.5 3745.9339334334336u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3755.708333833834u,0 3755.709333833834u,1.5 3758.6409539539536u,1.5 3758.641953953954u,0 3759.618493993994u,0 3759.619493993994u,1.5 3760.596034034034u,1.5 3760.597034034034u,0 3762.5511141141137u,0 3762.552114114114u,1.5 3764.506194194194u,1.5 3764.507194194194u,0 3766.461274274274u,0 3766.462274274274u,1.5 3770.3714344344344u,1.5 3770.3724344344346u,0 3775.259134634635u,0 3775.260134634635u,1.5 3776.2366746746743u,1.5 3776.2376746746745u,0 3778.1917547547546u,0 3778.192754754755u,1.5 3780.146834834835u,1.5 3780.147834834835u,0 3786.012075075075u,0 3786.013075075075u,1.5 3786.9896151151147u,1.5 3786.990615115115u,0 3787.967155155155u,0 3787.9681551551553u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3795.7874754754753u,0 3795.7884754754755u,1.5 3796.765015515515u,1.5 3796.7660155155154u,0 3797.7425555555556u,0 3797.7435555555558u,1.5 3799.697635635636u,1.5 3799.698635635636u,0 3801.6527157157157u,0 3801.653715715716u,1.5 3804.585335835836u,1.5 3804.586335835836u,0 3809.473036036036u,0 3809.474036036036u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3820.2259764764763u,0 3820.2269764764765u,1.5 3821.203516516516u,1.5 3821.2045165165164u,0 3822.1810565565565u,0 3822.1820565565567u,1.5 3829.023836836837u,1.5 3829.024836836837u,0 3830.9789169169167u,0 3830.979916916917u,1.5 3831.9564569569566u,1.5 3831.957456956957u,0 3833.911537037037u,0 3833.912537037037u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3839.776777277277u,0 3839.777777277277u,1.5 3840.754317317317u,1.5 3840.7553173173173u,0 3844.6644774774772u,0 3844.6654774774775u,1.5 3846.6195575575575u,1.5 3846.6205575575577u,0 3847.5970975975974u,0 3847.5980975975976u,1.5 3851.5072577577575u,1.5 3851.5082577577577u,0 3854.4398778778777u,0 3854.440877877878u,1.5 3855.4174179179176u,1.5 3855.418417917918u,0 3856.394957957958u,0 3856.395957957958u,1.5 3857.372497997998u,1.5 3857.373497997998u,0 3858.350038038038u,0 3858.351038038038u,1.5 3862.260198198198u,1.5 3862.261198198198u,0 3864.2152782782778u,0 3864.216278278278u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3870.080518518518u,0 3870.0815185185184u,1.5 3872.0355985985984u,1.5 3872.0365985985986u,0 3873.9906786786783u,0 3873.9916786786785u,1.5 3877.900838838839u,1.5 3877.901838838839u,0 3878.878378878879u,0 3878.8793788788794u,1.5 3879.8559189189186u,1.5 3879.856918918919u,0 3886.698699199199u,0 3886.699699199199u,1.5 3887.6762392392393u,1.5 3887.6772392392395u,0 3890.608859359359u,0 3890.6098593593592u,1.5 3892.5639394394393u,1.5 3892.5649394394395u,0 3903.31687987988u,0 3903.3178798798804u,1.5 3904.2944199199196u,1.5 3904.29541991992u,0 3905.27195995996u,0 3905.27295995996u,1.5 3907.22704004004u,1.5 3907.22804004004u,0 3908.20458008008u,0 3908.2055800800804u,1.5 3909.1821201201196u,1.5 3909.18312012012u,0 3910.1596601601605u,0 3910.1606601601607u,1.5 3913.09228028028u,1.5 3913.0932802802804u,0 3920.9126006006004u,0 3920.9136006006006u,1.5 3923.8452207207206u,1.5 3923.846220720721u,0 3924.822760760761u,0 3924.823760760761u,1.5 3928.7329209209206u,1.5 3928.733920920921u,0 3930.688001001001u,0 3930.689001001001u,1.5 3931.665541041041u,1.5 3931.666541041041u,0 3932.643081081081u,0 3932.6440810810814u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3937.530781281281u,1.5 3937.5317812812814u,0 3943.396021521521u,0 3943.3970215215213u,1.5 3944.373561561562u,1.5 3944.374561561562u,0 3947.3061816816817u,0 3947.307181681682u,1.5 3949.261261761762u,1.5 3949.262261761762u,0 3951.2163418418413u,0 3951.2173418418415u,1.5 3953.1714219219216u,1.5 3953.172421921922u,0 3954.1489619619624u,0 3954.1499619619626u,1.5 3955.126502002002u,1.5 3955.127502002002u,0 3956.104042042042u,0 3956.105042042042u,1.5 3957.081582082082u,1.5 3957.0825820820824u,0 3959.0366621621624u,0 3959.0376621621626u,1.5 3960.991742242242u,1.5 3960.992742242242u,0 3961.969282282282u,0 3961.9702822822824u,1.5 3964.9019024024024u,1.5 3964.9029024024026u,0 3965.879442442442u,0 3965.880442442442u,1.5 3966.8569824824826u,1.5 3966.857982482483u,0 3969.7896026026024u,0 3969.7906026026026u,1.5 3970.7671426426423u,1.5 3970.7681426426425u,0 3971.7446826826827u,0 3971.745682682683u,1.5 3972.7222227227226u,1.5 3972.7232227227228u,0 3974.677302802803u,0 3974.678302802803u,1.5 3976.632382882883u,1.5 3976.6333828828833u,0 3977.6099229229226u,0 3977.610922922923u,1.5 3978.5874629629634u,1.5 3978.5884629629636u,0 3985.430243243243u,0 3985.431243243243u,1.5 3986.407783283283u,1.5 3986.4087832832834u,0 3990.317943443443u,0 3990.318943443443u,1.5 3992.273023523523u,1.5 3992.2740235235233u,0 3994.2281036036034u,0 3994.2291036036036u,1.5 3995.2056436436433u,1.5 3995.2066436436435u,0 3996.1831836836836u,0 3996.184183683684u,1.5 3997.1607237237235u,1.5 3997.1617237237238u,0 3998.138263763764u,0 3998.139263763764u,1.5 4000.0933438438433u,1.5 4000.0943438438435u,0 4003.0259639639644u,0 4003.0269639639646u,1.5 4004.003504004004u,1.5 4004.004504004004u,0 4004.9810440440438u,0 4004.982044044044u,1.5 4005.958584084084u,1.5 4005.9595840840843u,0 4010.846284284284u,0 4010.8472842842843u,1.5 4013.7789044044043u,1.5 4013.7799044044045u,0 4018.6666046046043u,0 4018.6676046046045u,1.5 4019.6441446446443u,1.5 4019.6451446446445u,0 4023.554304804805u,0 4023.555304804805u,1.5 4024.5318448448443u,1.5 4024.5328448448445u,0 4025.509384884885u,0 4025.5103848848853u,1.5 4026.4869249249246u,1.5 4026.4879249249248u,0 4027.4644649649654u,0 4027.4654649649656u,1.5 4028.442005005005u,1.5 4028.443005005005u,0 4029.4195450450447u,0 4029.420545045045u,1.5 4031.374625125125u,1.5 4031.375625125125u,0 4032.3521651651654u,0 4032.3531651651656u,1.5 4033.329705205205u,1.5 4033.330705205205u,0 4035.284785285285u,0 4035.2857852852853u,1.5 4038.2174054054053u,1.5 4038.2184054054055u,0 4039.194945445445u,0 4039.195945445445u,1.5 4042.127565565566u,1.5 4042.128565565566u,0 4043.1051056056053u,0 4043.1061056056055u,1.5 4045.0601856856856u,1.5 4045.061185685686u,0 4046.0377257257255u,0 4046.0387257257257u,1.5 4047.992805805806u,1.5 4047.993805805806u,0 4048.9703458458453u,0 4048.9713458458455u,1.5 4049.947885885886u,1.5 4049.9488858858863u,0 4050.9254259259255u,0 4050.9264259259257u,1.5 4051.9029659659664u,1.5 4051.9039659659666u,0 4054.835586086086u,0 4054.8365860860863u,1.5 4055.813126126126u,1.5 4055.814126126126u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4072.431306806807u,0 4072.432306806807u,1.5 4075.3639269269265u,1.5 4075.3649269269267u,0 4077.319007007007u,0 4077.320007007007u,1.5 4080.251627127127u,1.5 4080.252627127127u,0 4081.2291671671674u,0 4081.2301671671676u,1.5 4083.1842472472467u,1.5 4083.185247247247u,0 4087.0944074074073u,0 4087.0954074074075u,1.5 4089.0494874874876u,1.5 4089.0504874874878u,0 4090.027027527527u,0 4090.0280275275272u,1.5 4093.9371876876876u,1.5 4093.938187687688u,0 4094.9147277277275u,0 4094.9157277277277u,1.5 4095.892267767768u,1.5 4095.893267767768u,0 4096.869807807808u,0 4096.870807807808u,1.5 4097.847347847847u,1.5 4097.848347847847u,0 4103.7125880880885u,0 4103.713588088089u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4106.645208208208u,0 4106.646208208208u,1.5 4111.532908408408u,1.5 4111.533908408408u,0 4112.510448448448u,0 4112.511448448448u,1.5 4113.487988488489u,1.5 4113.488988488489u,0 4120.330768768769u,0 4120.3317687687695u,1.5 4121.308308808809u,1.5 4121.309308808809u,0 4122.285848848848u,0 4122.286848848848u,1.5 4124.240928928929u,1.5 4124.241928928929u,0 4125.218468968969u,0 4125.2194689689695u,1.5 4129.128629129129u,1.5 4129.129629129129u,0 4130.106169169169u,0 4130.1071691691695u,1.5 4132.061249249249u,1.5 4132.062249249249u,0 4136.948949449449u,0 4136.949949449449u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4139.881569569569u,0 4139.88256956957u,1.5 4142.81418968969u,1.5 4142.81518968969u,0 4148.67942992993u,0 4148.68042992993u,1.5 4149.65696996997u,1.5 4149.6579699699705u,0 4150.63451001001u,0 4150.63551001001u,1.5 4154.54467017017u,1.5 4154.5456701701705u,0 4156.49975025025u,0 4156.50075025025u,1.5 4157.4772902902905u,1.5 4157.478290290291u,0 4160.40991041041u,0 4160.41091041041u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4162.3649904904905u,0 4162.365990490491u,1.5 4164.32007057057u,1.5 4164.321070570571u,0 4165.297610610611u,0 4165.298610610611u,1.5 4166.27515065065u,1.5 4166.27615065065u,0 4167.2526906906905u,0 4167.253690690691u,1.5 4168.23023073073u,1.5 4168.23123073073u,0 4172.140390890891u,0 4172.141390890891u,1.5 4178.005631131131u,1.5 4178.006631131131u,0 4178.983171171171u,0 4178.9841711711715u,1.5 4180.938251251251u,1.5 4180.939251251251u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4188.758571571571u,0 4188.7595715715715u,1.5 4191.6911916916915u,1.5 4191.692191691692u,0 4192.668731731731u,0 4192.669731731731u,1.5 4194.623811811812u,1.5 4194.624811811812u,0 4197.556431931932u,0 4197.557431931932u,1.5 4198.533971971972u,1.5 4198.5349719719725u,0 4199.511512012012u,0 4199.512512012012u,1.5 4200.489052052051u,1.5 4200.490052052051u,0 4201.4665920920925u,0 4201.467592092093u,1.5 4202.444132132132u,1.5 4202.445132132132u,0 4206.3542922922925u,0 4206.355292292293u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4210.264452452452u,1.5 4210.265452452452u,0 4212.219532532532u,0 4212.220532532532u,1.5 4213.197072572572u,1.5 4213.1980725725725u,0 4214.174612612613u,0 4214.175612612613u,1.5 4215.152152652652u,1.5 4215.153152652652u,0 4217.107232732732u,0 4217.108232732732u,1.5 4218.084772772773u,1.5 4218.085772772773u,0 4219.062312812813u,0 4219.063312812813u,1.5 4224.927553053052u,1.5 4224.928553053052u,0 4228.837713213213u,0 4228.838713213213u,1.5 4230.7927932932935u,1.5 4230.793793293294u,0 4231.770333333333u,0 4231.771333333333u,1.5 4234.702953453453u,1.5 4234.703953453453u,0 4236.658033533533u,0 4236.659033533533u,1.5 4238.613113613614u,1.5 4238.614113613614u,0 4240.5681936936935u,0 4240.569193693694u,1.5 4242.523273773774u,1.5 4242.524273773774u,0 4246.433433933934u,0 4246.434433933934u,1.5 4247.410973973974u,1.5 4247.411973973974u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4255.2312942942945u,1.5 4255.232294294295u,0 4256.208834334334u,0 4256.209834334334u,1.5 4257.186374374374u,1.5 4257.1873743743745u,0 4261.096534534534u,0 4261.097534534534u,1.5 4263.051614614615u,1.5 4263.052614614615u,0 4264.029154654655u,0 4264.030154654655u,1.5 4265.984234734734u,1.5 4265.985234734734u,0 4266.961774774775u,0 4266.962774774775u,1.5 4267.939314814815u,1.5 4267.940314814815u,0 4271.849474974975u,0 4271.850474974975u,1.5 4275.759635135135u,1.5 4275.760635135135u,0 4277.714715215215u,0 4277.715715215215u,1.5 4278.692255255256u,1.5 4278.693255255256u,0 4279.669795295295u,0 4279.670795295296u,1.5 4280.647335335335u,1.5 4280.648335335335u,0 4281.624875375375u,0 4281.6258753753755u,1.5 4284.5574954954955u,1.5 4284.558495495496u,0 4285.535035535535u,0 4285.536035535535u,1.5 4287.490115615616u,1.5 4287.491115615616u,0 4293.355355855856u,0 4293.356355855856u,1.5 4299.220596096096u,1.5 4299.221596096097u,0 4301.175676176176u,0 4301.176676176176u,1.5 4302.153216216216u,1.5 4302.154216216216u,0 4303.130756256257u,0 4303.131756256257u,1.5 4308.995996496496u,1.5 4308.996996496497u,0 4309.973536536536u,0 4309.974536536536u,1.5 4310.951076576576u,1.5 4310.9520765765765u,0 4315.838776776777u,0 4315.839776776777u,1.5 4316.816316816817u,1.5 4316.817316816817u,0 4317.793856856857u,0 4317.794856856857u,1.5 4318.7713968968965u,1.5 4318.772396896897u,0 4319.748936936937u,0 4319.749936936937u,1.5 4320.726476976977u,1.5 4320.727476976977u,0 4321.704017017017u,0 4321.705017017017u,1.5 4322.681557057057u,1.5 4322.682557057057u,0 4325.614177177177u,0 4325.615177177177u,1.5 4326.591717217217u,1.5 4326.592717217217u,0 4327.569257257258u,0 4327.570257257258u,1.5 4328.546797297297u,1.5 4328.547797297298u,0 4329.524337337337u,0 4329.525337337337u,1.5 4330.501877377377u,1.5 4330.502877377377u,0 4333.434497497497u,0 4333.435497497498u,1.5 4335.389577577577u,1.5 4335.3905775775775u,0 4338.322197697697u,0 4338.323197697698u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4342.232357857858u,1.5 4342.233357857858u,0 4344.187437937938u,0 4344.188437937938u,1.5 4345.164977977978u,1.5 4345.165977977978u,0 4351.030218218218u,0 4351.031218218218u,1.5 4352.007758258259u,1.5 4352.008758258259u,0 4352.985298298298u,0 4352.986298298299u,1.5 4353.962838338338u,1.5 4353.963838338338u,0 4354.940378378378u,0 4354.941378378378u,1.5 4357.872998498498u,1.5 4357.873998498499u,0 4358.850538538538u,0 4358.851538538538u,1.5 4359.828078578578u,1.5 4359.829078578578u,0 4360.805618618619u,0 4360.806618618619u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4371.558559059059u,1.5 4371.559559059059u,0 4374.491179179179u,0 4374.492179179179u,1.5 4375.468719219219u,1.5 4375.469719219219u,0 4376.44625925926u,0 4376.44725925926u,1.5 4377.423799299299u,1.5 4377.4247992993u,0 4379.378879379379u,0 4379.379879379379u,1.5 4384.266579579579u,1.5 4384.267579579579u,0 4387.199199699699u,0 4387.2001996997u,1.5 4388.176739739739u,1.5 4388.177739739739u,0 4389.15427977978u,0 4389.15527977978u,1.5 4390.13181981982u,1.5 4390.13281981982u,0 4392.086899899899u,0 4392.0878998999u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.01952002002u,1.5 4395.02052002002u,0 4397.95214014014u,0 4397.95314014014u,1.5 4402.83984034034u,1.5 4402.84084034034u,0 4403.81738038038u,0 4403.81838038038u,1.5 4405.772460460461u,1.5 4405.773460460461u,0 4407.72754054054u,0 4407.72854054054u,1.5 4408.70508058058u,1.5 4408.70608058058u,0 4409.682620620621u,0 4409.683620620621u,1.5 4410.660160660661u,1.5 4410.661160660661u,0 4412.61524074074u,0 4412.61624074074u,1.5 4414.570320820821u,1.5 4414.571320820821u,0 4415.547860860861u,0 4415.548860860861u,1.5 4417.502940940941u,1.5 4417.503940940941u,0 4418.480480980981u,0 4418.481480980981u,1.5 4422.390641141141u,1.5 4422.391641141141u,0 4424.345721221221u,0 4424.346721221221u,1.5 4425.323261261262u,1.5 4425.324261261262u,0 4426.300801301301u,0 4426.301801301302u,1.5 4427.278341341341u,1.5 4427.279341341341u,0 4430.210961461462u,0 4430.211961461462u,1.5 4431.188501501501u,1.5 4431.189501501502u,0 4432.166041541541u,0 4432.167041541541u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4439.008821821822u,1.5 4439.009821821822u,0 4441.941441941942u,0 4441.942441941942u,1.5 4443.896522022022u,1.5 4443.897522022022u,0 4444.874062062062u,0 4444.875062062062u,1.5 4446.829142142142u,1.5 4446.830142142142u,0 4448.784222222222u,0 4448.785222222222u,1.5 4449.761762262263u,1.5 4449.762762262263u,0 4450.739302302302u,0 4450.740302302303u,1.5 4451.716842342342u,1.5 4451.717842342342u,0 4453.6719224224225u,0 4453.672922422423u,1.5 4454.649462462463u,1.5 4454.650462462463u,0 4456.604542542542u,0 4456.605542542542u,1.5 4460.514702702702u,1.5 4460.515702702703u,0 4467.357482982983u,0 4467.358482982983u,1.5 4468.335023023023u,1.5 4468.336023023023u,0 4469.312563063063u,0 4469.313563063063u,1.5 4471.267643143143u,1.5 4471.268643143143u,0 4472.245183183183u,0 4472.246183183183u,1.5 4473.222723223223u,1.5 4473.223723223223u,0 4474.200263263264u,0 4474.201263263264u,1.5 4475.177803303303u,1.5 4475.1788033033035u,0 4476.155343343343u,0 4476.156343343343u,1.5 4478.1104234234235u,1.5 4478.111423423424u,0 4479.087963463464u,0 4479.088963463464u,1.5 4482.9981236236235u,1.5 4482.999123623624u,0 4485.930743743743u,0 4485.931743743743u,1.5 4491.795983983984u,1.5 4491.796983983984u,0 4492.773524024024u,0 4492.774524024024u,1.5 4494.728604104104u,1.5 4494.7296041041045u,0 4496.683684184184u,0 4496.684684184184u,1.5 4503.526464464465u,1.5 4503.527464464465u,0 4504.504004504504u,0 4504.5050045045045u,1.5 4505.481544544544u,1.5 4505.482544544544u,0 4508.414164664665u,0 4508.415164664665u,1.5 4510.369244744744u,1.5 4510.370244744744u,0 4511.346784784785u,0 4511.347784784785u,1.5 4514.279404904904u,1.5 4514.280404904905u,0 4515.256944944945u,0 4515.257944944945u,1.5 4519.167105105105u,1.5 4519.1681051051055u,0 4520.144645145145u,0 4520.145645145145u,1.5 4522.099725225225u,1.5 4522.100725225225u,0 4523.077265265266u,0 4523.078265265266u,1.5 4525.032345345345u,1.5 4525.033345345345u,0 4526.9874254254255u,0 4526.988425425426u,1.5 4528.942505505505u,1.5 4528.9435055055055u,0 4529.920045545545u,0 4529.921045545545u,1.5 4531.8751256256255u,1.5 4531.876125625626u,0 4536.7628258258255u,0 4536.763825825826u,1.5 4537.740365865866u,1.5 4537.741365865866u,0 4539.695445945946u,0 4539.696445945946u,1.5 4540.672985985986u,1.5 4540.673985985986u,0 4541.650526026026u,0 4541.651526026026u,1.5 4544.583146146146u,1.5 4544.584146146146u,0 4545.560686186186u,0 4545.561686186186u,1.5 4546.538226226226u,1.5 4546.539226226226u,0 4548.493306306306u,0 4548.4943063063065u,1.5 4550.448386386386u,1.5 4550.449386386386u,0 4551.4259264264265u,0 4551.426926426427u,1.5 4555.336086586587u,1.5 4555.337086586587u,0 4556.3136266266265u,0 4556.314626626627u,1.5 4562.178866866867u,1.5 4562.179866866867u,0 4563.156406906906u,0 4563.1574069069065u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4569.021647147147u,0 4569.022647147147u,1.5 4569.999187187187u,1.5 4570.000187187187u,0 4576.841967467468u,0 4576.842967467468u,1.5 4577.819507507507u,1.5 4577.8205075075075u,0 4578.797047547547u,0 4578.798047547547u,1.5 4583.684747747748u,1.5 4583.685747747748u,0 4585.6398278278275u,0 4585.640827827828u,1.5 4586.617367867868u,1.5 4586.618367867868u,0 4587.594907907907u,0 4587.5959079079075u,1.5 4588.572447947948u,1.5 4588.573447947948u,0 4590.5275280280275u,0 4590.528528028028u,1.5 4591.505068068068u,1.5 4591.506068068068u,0 4597.370308308308u,0 4597.3713083083085u,1.5 4600.3029284284285u,1.5 4600.303928428429u,0 4601.280468468469u,0 4601.281468468469u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4607.145708708708u,0 4607.1467087087085u,1.5 4608.123248748749u,1.5 4608.124248748749u,0 4613.988488988989u,0 4613.989488988989u,1.5 4614.9660290290285u,1.5 4614.967029029029u,0 4615.943569069069u,0 4615.944569069069u,1.5 4616.921109109109u,1.5 4616.922109109109u,0 4617.898649149149u,0 4617.899649149149u,1.5 4620.83126926927u,1.5 4620.83226926927u,0 4622.786349349349u,0 4622.787349349349u,1.5 4623.763889389389u,1.5 4623.764889389389u,0 4627.674049549549u,0 4627.675049549549u,1.5 4629.6291296296295u,1.5 4629.63012962963u,0 4630.60666966967u,0 4630.60766966967u,1.5 4633.53928978979u,1.5 4633.54028978979u,0 4635.49436986987u,0 4635.49536986987u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4640.38207007007u,0 4640.38307007007u,1.5 4641.35961011011u,1.5 4641.36061011011u,0 4643.31469019019u,0 4643.31569019019u,1.5 4645.269770270271u,1.5 4645.270770270271u,0 4646.24731031031u,0 4646.24831031031u,1.5 4649.17993043043u,1.5 4649.180930430431u,0 4651.13501051051u,0 4651.1360105105105u,1.5 4652.11255055055u,1.5 4652.11355055055u,0 4653.090090590591u,0 4653.091090590591u,1.5 4654.06763063063u,1.5 4654.068630630631u,0 4655.045170670671u,0 4655.046170670671u,1.5 4657.000250750751u,1.5 4657.001250750751u,0 4657.977790790791u,0 4657.978790790791u,1.5 4658.9553308308305u,1.5 4658.956330830831u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4665.798111111111u,0 4665.799111111111u,1.5 4669.708271271272u,1.5 4669.709271271272u,0 4670.685811311311u,0 4670.686811311311u,1.5 4671.663351351351u,1.5 4671.664351351351u,0 4680.461211711711u,0 4680.4622117117115u,1.5 4682.416291791792u,1.5 4682.417291791792u,0 4683.393831831831u,0 4683.394831831832u,1.5 4685.348911911911u,1.5 4685.3499119119115u,0 4686.326451951952u,0 4686.327451951952u,1.5 4687.303991991992u,1.5 4687.304991991992u,0 4688.2815320320315u,0 4688.282532032032u,1.5 4689.259072072072u,1.5 4689.260072072072u,0 4691.214152152152u,0 4691.215152152152u,1.5 4692.191692192192u,1.5 4692.192692192192u,0 4693.1692322322315u,0 4693.170232232232u,1.5 4697.079392392392u,1.5 4697.080392392392u,0 4698.056932432432u,0 4698.057932432433u,1.5 4699.034472472473u,1.5 4699.035472472473u,0 4700.012012512512u,0 4700.013012512512u,1.5 4700.989552552552u,1.5 4700.990552552552u,0 4702.944632632632u,0 4702.945632632633u,1.5 4704.899712712712u,1.5 4704.900712712712u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4709.787412912912u,1.5 4709.7884129129125u,0 4713.697573073073u,0 4713.698573073073u,1.5 4718.585273273274u,1.5 4718.586273273274u,0 4720.540353353353u,0 4720.541353353353u,1.5 4722.495433433433u,1.5 4722.496433433434u,0 4725.428053553553u,0 4725.429053553553u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4734.225913913913u,0 4734.226913913913u,1.5 4735.203453953954u,1.5 4735.204453953954u,0 4736.180993993994u,0 4736.181993993994u,1.5 4740.091154154154u,1.5 4740.092154154154u,0 4744.001314314314u,0 4744.002314314314u,1.5 4744.978854354354u,1.5 4744.979854354354u,0 4745.956394394394u,0 4745.957394394394u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4753.776714714714u,0 4753.777714714714u,1.5 4754.7542547547555u,1.5 4754.755254754756u,0 4755.731794794795u,0 4755.732794794795u,1.5 4756.709334834834u,1.5 4756.710334834835u,0 4757.686874874875u,0 4757.687874874875u,1.5 4760.619494994995u,1.5 4760.620494994995u,0 4761.597035035034u,0 4761.598035035035u,1.5 4763.552115115115u,1.5 4763.553115115115u,0 4767.462275275276u,0 4767.463275275276u,1.5 4770.394895395395u,1.5 4770.395895395395u,0 4772.349975475476u,0 4772.350975475476u,1.5 4774.305055555556u,1.5 4774.306055555556u,0 4778.215215715715u,0 4778.216215715715u,1.5 4781.147835835835u,1.5 4781.148835835836u,0 4784.0804559559565u,0 4784.081455955957u,1.5 4786.035536036035u,1.5 4786.036536036036u,0 4787.990616116116u,0 4787.991616116116u,1.5 4792.878316316316u,1.5 4792.879316316316u,0 4794.833396396396u,0 4794.834396396396u,1.5 4797.766016516516u,1.5 4797.767016516516u,0 4799.721096596597u,0 4799.722096596597u,1.5 4804.608796796797u,1.5 4804.609796796797u,0 4809.496496996997u,0 4809.497496996997u,1.5 4810.474037037036u,1.5 4810.475037037037u,0 4811.451577077077u,0 4811.452577077077u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4816.339277277278u,0 4816.340277277278u,1.5 4817.316817317317u,1.5 4817.317817317317u,0 4819.271897397397u,0 4819.272897397397u,1.5 4822.204517517517u,1.5 4822.205517517517u,0 4824.159597597598u,0 4824.160597597598u,1.5 4825.137137637637u,1.5 4825.138137637638u,0 4826.114677677678u,0 4826.115677677678u,1.5 4827.092217717717u,1.5 4827.093217717717u,0 4831.002377877878u,0 4831.003377877878u,1.5 4831.979917917918u,1.5 4831.980917917918u,0 4832.9574579579585u,0 4832.958457957959u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4843.710398398398u,0 4843.711398398398u,1.5 4844.687938438438u,1.5 4844.6889384384385u,0 4845.665478478479u,0 4845.666478478479u,1.5 4849.575638638638u,1.5 4849.5766386386385u,0 4850.553178678679u,0 4850.554178678679u,1.5 4851.530718718718u,1.5 4851.531718718718u,0 4852.508258758759u,0 4852.50925875876u,1.5 4853.485798798799u,1.5 4853.486798798799u,0 4854.463338838838u,0 4854.464338838839u,1.5 4855.440878878879u,1.5 4855.441878878879u,0 4857.395958958959u,0 4857.39695895896u,1.5 4865.21627927928u,1.5 4865.21727927928u,0 4870.10397947948u,0 4870.10497947948u,1.5 4872.0590595595595u,1.5 4872.06005955956u,0 4873.0365995996u,0 4873.0375995996u,1.5 4876.94675975976u,1.5 4876.947759759761u,0 4877.9242997998u,0 4877.9252997998u,1.5 4878.901839839839u,1.5 4878.9028398398395u,0 4879.87937987988u,0 4879.88037987988u,1.5 4880.85691991992u,1.5 4880.85791991992u,0 4881.83445995996u,0 4881.835459959961u,1.5 4885.74462012012u,1.5 4885.74562012012u,0 4886.7221601601605u,0 4886.723160160161u,1.5 4890.63232032032u,1.5 4890.63332032032u,0 4891.6098603603605u,0 4891.610860360361u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4895.52002052052u,0 4895.52102052052u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4903.34034084084u,0 4903.3413408408405u,1.5 4905.295420920921u,1.5 4905.296420920921u,0 4906.272960960961u,0 4906.273960960962u,1.5 4907.250501001001u,1.5 4907.251501001001u,0 4908.22804104104u,0 4908.229041041041u,1.5 4911.160661161161u,1.5 4911.161661161162u,0 4912.138201201201u,0 4912.139201201201u,1.5 4914.093281281282u,1.5 4914.094281281282u,0 4917.025901401401u,0 4917.026901401401u,1.5 4918.980981481482u,1.5 4918.981981481482u,0 4919.958521521521u,0 4919.959521521521u,1.5 4920.9360615615615u,1.5 4920.937061561562u,0 4921.913601601602u,0 4921.914601601602u,1.5 4923.868681681682u,1.5 4923.869681681682u,0 4924.846221721721u,0 4924.847221721721u,1.5 4930.711461961962u,1.5 4930.712461961963u,0 4931.689002002002u,0 4931.690002002002u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4935.599162162162u,1.5 4935.600162162163u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4939.509322322322u,0 4939.510322322322u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 4945.3745625625625u,0 4945.375562562563u,1.5 4946.352102602603u,1.5 4946.353102602603u,0 4950.262262762763u,0 4950.263262762764u,1.5 4956.127503003003u,1.5 4956.128503003003u,0 4957.105043043042u,0 4957.1060430430425u,1.5 4964.925363363363u,1.5 4964.926363363364u,0 4965.902903403403u,0 4965.903903403403u,1.5 4969.813063563563u,1.5 4969.814063563564u,0 4970.790603603604u,0 4970.791603603604u,1.5 4971.768143643643u,1.5 4971.7691436436435u,0 4972.745683683684u,0 4972.746683683684u,1.5 4973.723223723723u,1.5 4973.724223723723u,0 4974.700763763764u,0 4974.701763763765u,1.5 4976.655843843843u,1.5 4976.6568438438435u,0 4977.633383883884u,0 4977.634383883884u,1.5 4978.610923923924u,1.5 4978.611923923924u,0 4983.498624124124u,0 4983.499624124124u,1.5 4984.476164164164u,1.5 4984.477164164165u,0 4985.453704204204u,0 4985.454704204204u,1.5 4986.431244244243u,1.5 4986.4322442442435u,0 4988.386324324324u,0 4988.387324324324u,1.5 4989.363864364364u,1.5 4989.364864364365u,0 4999.139264764765u,0 4999.140264764766u,1.5 5000.116804804805u,1.5 5000.117804804805u,0 5003.049424924925u,0 5003.050424924925u,1.5 5005.004505005005u,1.5 5005.005505005005u,0 5005.982045045044u,0 5005.9830450450445u,1.5 5007.937125125125u,1.5 5007.938125125125u,0 5014.779905405405u,0 5014.780905405405u,1.5 5016.734985485486u,1.5 5016.735985485486u,0 5017.712525525525u,0 5017.713525525525u,1.5 5018.690065565565u,1.5 5018.691065565566u,0 5020.645145645645u,0 5020.646145645645u,1.5 5024.555305805806u,1.5 5024.556305805806u,0 5025.532845845845u,0 5025.5338458458455u,1.5 5026.510385885886u,1.5 5026.511385885886u,0 5028.465465965966u,0 5028.466465965967u,1.5 5029.443006006006u,1.5 5029.444006006006u,0 5031.398086086087u,0 5031.399086086087u,1.5 5033.353166166166u,1.5 5033.354166166167u,0 5034.330706206206u,0 5034.331706206206u,1.5 5042.151026526526u,1.5 5042.152026526526u,0 5043.128566566566u,0 5043.129566566567u,1.5 5044.106106606607u,1.5 5044.107106606607u,0 5045.083646646646u,0 5045.084646646646u,1.5 5048.993806806807u,1.5 5048.994806806807u,0 5049.971346846846u,0 5049.972346846846u,1.5 5050.948886886887u,1.5 5050.949886886887u,0 5052.903966966967u,0 5052.904966966968u,1.5 5053.881507007007u,1.5 5053.882507007007u,0 5054.859047047046u,0 5054.8600470470465u,1.5 5057.791667167167u,1.5 5057.792667167168u,0 5059.746747247247u,0 5059.747747247247u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5067.567067567567u,1.5 5067.568067567568u,0 5068.544607607608u,0 5068.545607607608u,1.5 5071.477227727727u,1.5 5071.478227727727u,0 5072.454767767768u,0 5072.4557677677685u,1.5 5074.409847847847u,1.5 5074.410847847847u,0 5075.387387887888u,0 5075.388387887888u,1.5 5077.342467967968u,1.5 5077.3434679679685u,0 5078.320008008008u,0 5078.321008008008u,1.5 5079.297548048047u,1.5 5079.298548048047u,0 5081.252628128128u,0 5081.253628128128u,1.5 5082.230168168168u,1.5 5082.231168168169u,0 5084.185248248248u,0 5084.186248248248u,1.5 5085.1627882882885u,1.5 5085.163788288289u,0 5087.117868368368u,0 5087.118868368369u,1.5 5088.095408408408u,1.5 5088.096408408408u,0 5089.072948448448u,0 5089.073948448448u,1.5 5092.983108608609u,1.5 5092.984108608609u,0 5103.736049049048u,0 5103.737049049048u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5108.623749249249u,0 5108.624749249249u,1.5 5113.511449449449u,1.5 5113.512449449449u,0 5116.444069569569u,0 5116.44506956957u,1.5 5118.399149649649u,1.5 5118.400149649649u,0 5121.33176976977u,0 5121.3327697697705u,1.5 5122.30930980981u,1.5 5122.31030980981u,0 5123.286849849849u,0 5123.287849849849u,1.5 5129.1520900900905u,1.5 5129.153090090091u,0 5131.10717017017u,0 5131.1081701701705u,1.5 5132.08471021021u,1.5 5132.08571021021u,0 5134.0397902902905u,0 5134.040790290291u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5138.9274904904905u,0 5138.928490490491u,1.5 5141.860110610611u,1.5 5141.861110610611u,0 5142.83765065065u,0 5142.83865065065u,1.5 5143.8151906906905u,1.5 5143.816190690691u,0 5148.702890890891u,0 5148.703890890891u,1.5 5154.568131131131u,1.5 5154.569131131131u,0 5155.545671171171u,0 5155.5466711711715u,1.5 5156.523211211211u,1.5 5156.524211211211u,0 5157.500751251251u,0 5157.501751251251u,1.5 5159.455831331331u,1.5 5159.456831331331u,0 5161.410911411411u,0 5161.411911411411u,1.5 5163.3659914914915u,1.5 5163.366991491492u,0 5164.343531531531u,0 5164.344531531531u,1.5 5167.276151651651u,1.5 5167.277151651651u,0 5169.231231731731u,0 5169.232231731731u,1.5 5170.208771771772u,1.5 5170.2097717717725u,0 5173.1413918918915u,0 5173.142391891892u,1.5 5174.118931931932u,1.5 5174.119931931932u,0 5175.096471971972u,0 5175.0974719719725u,1.5 5180.961712212212u,1.5 5180.962712212212u,0 5181.939252252252u,0 5181.940252252252u,1.5 5182.9167922922925u,1.5 5182.917792292293u,0 5185.849412412412u,0 5185.850412412412u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5187.8044924924925u,0 5187.805492492493u,1.5 5189.759572572572u,1.5 5189.7605725725725u,0 5190.737112612613u,0 5190.738112612613u,1.5 5191.714652652652u,1.5 5191.715652652652u,0 5193.669732732732u,0 5193.670732732732u,1.5 5194.647272772773u,1.5 5194.648272772773u,0 5197.5798928928925u,0 5197.580892892893u,1.5 5203.445133133133u,1.5 5203.446133133133u,0 5207.3552932932935u,0 5207.356293293294u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5211.265453453453u,0 5211.266453453453u,1.5 5213.220533533533u,1.5 5213.221533533533u,0 5214.198073573573u,0 5214.1990735735735u,1.5 5216.153153653653u,1.5 5216.154153653653u,0 5217.1306936936935u,0 5217.131693693694u,1.5 5218.108233733733u,1.5 5218.109233733733u,0 5219.085773773774u,0 5219.086773773774u,1.5 5220.063313813814u,1.5 5220.064313813814u,0 5221.040853853853u,0 5221.041853853853u,1.5 5223.973473973974u,1.5 5223.974473973974u,0 5224.951014014014u,0 5224.952014014014u,1.5 5225.928554054053u,1.5 5225.929554054053u,0 5228.861174174174u,0 5228.8621741741745u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5235.703954454454u,1.5 5235.704954454454u,0 5239.614114614615u,0 5239.615114614615u,1.5 5244.501814814815u,1.5 5244.502814814815u,0 5245.479354854854u,0 5245.480354854854u,1.5 5246.4568948948945u,1.5 5246.457894894895u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5258.187375375375u,1.5 5258.1883753753755u,0 5259.164915415415u,0 5259.165915415415u,1.5 5261.1199954954955u,1.5 5261.120995495496u,0 5262.097535535535u,0 5262.098535535535u,1.5 5263.075075575575u,1.5 5263.0760755755755u,0 5266.0076956956955u,0 5266.008695695696u,1.5 5266.985235735735u,1.5 5266.986235735735u,0 5271.872935935936u,0 5271.873935935936u,1.5 5274.805556056056u,1.5 5274.806556056056u,0 5281.648336336336u,0 5281.649336336336u,1.5 5282.625876376376u,1.5 5282.6268763763765u,0 5284.580956456457u,0 5284.581956456457u,1.5 5288.491116616617u,1.5 5288.492116616617u,0 5292.401276776777u,0 5292.402276776777u,1.5 5297.288976976977u,1.5 5297.289976976977u,0 5300.221597097097u,0 5300.222597097098u,1.5 5301.199137137137u,1.5 5301.200137137137u,0 5303.154217217217u,0 5303.155217217217u,1.5 5309.019457457458u,1.5 5309.020457457458u,0 5310.974537537537u,0 5310.975537537537u,1.5 5311.952077577577u,1.5 5311.9530775775775u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5316.839777777778u,0 5316.840777777778u,1.5 5319.7723978978975u,1.5 5319.773397897898u,0 5327.592718218218u,0 5327.593718218218u,1.5 5331.502878378378u,1.5 5331.503878378378u,0 5332.480418418419u,0 5332.481418418419u,1.5 5333.457958458459u,1.5 5333.458958458459u,0 5339.323198698698u,0 5339.324198698699u,1.5 5344.210898898898u,1.5 5344.211898898899u,0 5345.188438938939u,0 5345.189438938939u,1.5 5347.143519019019u,1.5 5347.144519019019u,0 5348.121059059059u,0 5348.122059059059u,1.5 5350.076139139139u,1.5 5350.077139139139u,0 5352.031219219219u,0 5352.032219219219u,1.5 5357.89645945946u,1.5 5357.89745945946u,0 5359.851539539539u,0 5359.852539539539u,1.5 5360.829079579579u,1.5 5360.830079579579u,0 5365.71677977978u,0 5365.71777977978u,1.5 5369.62693993994u,1.5 5369.62793993994u,0 5370.60447997998u,0 5370.60547997998u,1.5 5371.58202002002u,1.5 5371.58302002002u,0 5376.46972022022u,0 5376.47072022022u,1.5 5377.447260260261u,1.5 5377.448260260261u,0 5378.4248003003u,0 5378.425800300301u,1.5 5380.37988038038u,1.5 5380.38088038038u,0 5382.334960460461u,0 5382.335960460461u,1.5 5387.222660660661u,1.5 5387.223660660661u,0 5392.110360860861u,0 5392.111360860861u,1.5 5393.0879009009u,1.5 5393.088900900901u,0 5396.020521021021u,0 5396.021521021021u,1.5 5400.908221221221u,1.5 5400.909221221221u,0 5401.885761261262u,0 5401.886761261262u,1.5 5404.818381381381u,1.5 5404.819381381381u,0 5408.728541541541u,0 5408.729541541541u,1.5 5409.706081581581u,1.5 5409.707081581581u,0 5411.661161661662u,0 5411.662161661662u,1.5 5412.638701701701u,1.5 5412.639701701702u,0 5415.571321821822u,0 5415.572321821822u,1.5 5417.526401901901u,1.5 5417.527401901902u,0 5418.503941941942u,0 5418.504941941942u,1.5 5421.436562062062u,1.5 5421.437562062062u,0 5422.414102102102u,0 5422.4151021021025u,1.5 5423.391642142142u,1.5 5423.392642142142u,0 5424.369182182182u,0 5424.370182182182u,1.5 5425.346722222222u,1.5 5425.347722222222u,0 5433.167042542542u,0 5433.168042542542u,1.5 5434.144582582582u,1.5 5434.145582582582u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5442.942442942943u,1.5 5442.943442942943u,0 5444.897523023023u,0 5444.898523023023u,1.5 5446.852603103103u,1.5 5446.8536031031035u,0 5447.830143143143u,0 5447.831143143143u,1.5 5448.807683183183u,1.5 5448.808683183183u,0 5450.762763263264u,0 5450.763763263264u,1.5 5452.717843343343u,1.5 5452.718843343343u,0 5456.628003503503u,0 5456.629003503504u,1.5 5458.583083583583u,1.5 5458.584083583583u,0 5459.5606236236235u,0 5459.561623623624u,1.5 5461.515703703703u,1.5 5461.516703703704u,0 5466.403403903903u,0 5466.404403903904u,1.5 5467.380943943944u,1.5 5467.381943943944u,0 5468.358483983984u,0 5468.359483983984u,1.5 5469.336024024024u,1.5 5469.337024024024u,0 5471.291104104104u,0 5471.2921041041045u,1.5 5473.246184184184u,1.5 5473.247184184184u,0 5474.223724224224u,0 5474.224724224224u,1.5 5475.201264264265u,1.5 5475.202264264265u,0 5476.178804304304u,0 5476.1798043043045u,1.5 5478.133884384384u,1.5 5478.134884384384u,0 5479.1114244244245u,0 5479.112424424425u,1.5 5481.066504504504u,1.5 5481.0675045045045u,0 5482.044044544544u,0 5482.045044544544u,1.5 5483.9991246246245u,1.5 5484.000124624625u,0 5484.976664664665u,0 5484.977664664665u,1.5 5490.841904904904u,1.5 5490.842904904905u,0 5491.819444944945u,0 5491.820444944945u,1.5 5492.796984984985u,1.5 5492.797984984985u,0 5495.729605105105u,0 5495.7306051051055u,1.5 5497.684685185185u,1.5 5497.685685185185u,0 5498.662225225225u,0 5498.663225225225u,1.5 5503.5499254254255u,1.5 5503.550925425426u,0 5504.527465465466u,0 5504.528465465466u,1.5 5511.370245745745u,1.5 5511.371245745745u,0 5513.3253258258255u,0 5513.326325825826u,1.5 5520.168106106106u,1.5 5520.1691061061065u,0 5522.123186186186u,0 5522.124186186186u,1.5 5524.078266266267u,1.5 5524.079266266267u,0 5525.055806306306u,0 5525.0568063063065u,1.5 5527.9884264264265u,1.5 5527.989426426427u,0 5528.965966466467u,0 5528.966966466467u,1.5 5529.943506506506u,1.5 5529.9445065065065u,0 5533.853666666667u,0 5533.854666666667u,1.5 5534.831206706706u,1.5 5534.8322067067065u,0 5539.718906906906u,0 5539.7199069069065u,1.5 5544.606607107107u,1.5 5544.6076071071075u,0 5547.539227227227u,0 5547.540227227227u,1.5 5548.516767267268u,1.5 5548.517767267268u,0 5551.449387387387u,0 5551.450387387387u,1.5 5553.404467467468u,1.5 5553.405467467468u,0 5554.382007507507u,0 5554.3830075075075u,1.5 5557.3146276276275u,1.5 5557.315627627628u,0 5559.269707707707u,0 5559.2707077077075u,1.5 5564.157407907907u,1.5 5564.1584079079075u,0 5568.067568068068u,0 5568.068568068068u,1.5 5569.045108108108u,1.5 5569.0461081081085u,0 5574.910348348348u,0 5574.911348348348u,1.5 5575.887888388388u,1.5 5575.888888388388u,0 5578.820508508508u,0 5578.8215085085085u,1.5 5584.685748748749u,1.5 5584.686748748749u,0 5585.663288788789u,0 5585.664288788789u,1.5 5587.618368868869u,1.5 5587.619368868869u,0 5596.4162292292285u,0 5596.417229229229u,1.5 5598.371309309309u,1.5 5598.3723093093095u,0 5600.326389389389u,0 5600.327389389389u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5602.28146946947u,0 5602.28246946947u,1.5 5604.236549549549u,1.5 5604.237549549549u,0 5606.1916296296295u,0 5606.19262962963u,1.5 5607.16916966967u,1.5 5607.17016966967u,0 5608.146709709709u,0 5608.1477097097095u,1.5 5609.12424974975u,1.5 5609.12524974975u,0 5614.01194994995u,0 5614.01294994995u,1.5 5614.98948998999u,1.5 5614.99048998999u,0 5615.9670300300295u,0 5615.96803003003u,1.5 5616.94457007007u,1.5 5616.94557007007u,0 5618.89965015015u,0 5618.90065015015u,1.5 5619.87719019019u,1.5 5619.87819019019u,0 5620.8547302302295u,0 5620.85573023023u,1.5 5623.78735035035u,1.5 5623.78835035035u,0 5626.719970470471u,0 5626.720970470471u,1.5 5627.69751051051u,1.5 5627.6985105105105u,0 5628.67505055055u,0 5628.67605055055u,1.5 5630.63013063063u,1.5 5630.631130630631u,0 5631.607670670671u,0 5631.608670670671u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5641.383071071071u,0 5641.384071071071u,1.5 5642.360611111111u,1.5 5642.361611111111u,0 5643.338151151151u,0 5643.339151151151u,1.5 5644.315691191191u,1.5 5644.316691191191u,0 5645.2932312312305u,0 5645.294231231231u,1.5 5647.248311311311u,1.5 5647.249311311311u,0 5650.180931431431u,0 5650.181931431432u,1.5 5652.136011511511u,1.5 5652.137011511511u,0 5656.046171671672u,0 5656.047171671672u,1.5 5657.023711711711u,1.5 5657.0247117117115u,0 5658.001251751752u,0 5658.002251751752u,1.5 5659.956331831831u,1.5 5659.957331831832u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5662.888951951952u,1.5 5662.889951951952u,0 5668.754192192192u,0 5668.755192192192u,1.5 5672.664352352352u,1.5 5672.665352352352u,0 5674.619432432432u,0 5674.620432432433u,1.5 5675.596972472473u,1.5 5675.597972472473u,0 5680.484672672673u,0 5680.485672672673u,1.5 5685.372372872873u,1.5 5685.373372872873u,0 5686.349912912912u,0 5686.3509129129125u,1.5 5687.327452952953u,1.5 5687.328452952953u,0 5692.215153153153u,0 5692.216153153153u,1.5 5693.192693193193u,1.5 5693.193693193193u,0 5694.1702332332325u,0 5694.171233233233u,1.5 5696.125313313313u,1.5 5696.126313313313u,0 5698.080393393393u,0 5698.081393393393u,1.5 5700.035473473474u,1.5 5700.036473473474u,0 5701.990553553553u,0 5701.991553553553u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5712.743493993994u,0 5712.744493993994u,1.5 5713.721034034033u,1.5 5713.722034034034u,0 5714.698574074074u,0 5714.699574074074u,1.5 5719.586274274275u,1.5 5719.587274274275u,0 5721.541354354354u,0 5721.542354354354u,1.5 5722.518894394394u,1.5 5722.519894394394u,0 5723.496434434434u,0 5723.497434434435u,1.5 5724.473974474475u,1.5 5724.474974474475u,0 5725.451514514514u,0 5725.452514514514u,1.5 5728.384134634634u,1.5 5728.385134634635u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5731.316754754755u,0 5731.317754754755u,1.5 5732.294294794795u,1.5 5732.295294794795u,0 5735.226914914914u,0 5735.227914914914u,1.5 5736.204454954955u,1.5 5736.205454954955u,0 5737.181994994995u,0 5737.182994994995u,1.5 5739.137075075075u,1.5 5739.138075075075u,0 5740.114615115115u,0 5740.115615115115u,1.5 5741.092155155155u,1.5 5741.093155155155u,0 5745.002315315315u,0 5745.003315315315u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5753.800175675676u,0 5753.801175675676u,1.5 5760.6429559559565u,1.5 5760.643955955957u,0 5762.598036036035u,0 5762.599036036036u,1.5 5763.575576076076u,1.5 5763.576576076076u,0 5766.508196196196u,0 5766.509196196196u,1.5 5767.485736236235u,1.5 5767.486736236236u,0 5768.463276276277u,0 5768.464276276277u,1.5 5769.440816316316u,1.5 5769.441816316316u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5775.3060565565565u,0 5775.307056556557u,1.5 5776.283596596597u,1.5 5776.284596596597u,0 5777.261136636636u,0 5777.262136636637u,1.5 5778.238676676677u,1.5 5778.239676676677u,0 5779.216216716716u,0 5779.217216716716u,1.5 5780.1937567567575u,1.5 5780.194756756758u,0 5781.171296796797u,0 5781.172296796797u,1.5 5782.148836836836u,1.5 5782.149836836837u,0 5785.0814569569575u,0 5785.082456956958u,1.5 5791.924237237236u,1.5 5791.925237237237u,0 5794.8568573573575u,0 5794.857857357358u,1.5 5795.834397397397u,1.5 5795.835397397397u,0 5796.811937437437u,0 5796.8129374374375u,1.5 5797.789477477478u,1.5 5797.790477477478u,0 5798.767017517517u,0 5798.768017517517u,1.5 5802.677177677678u,1.5 5802.678177677678u,0 5803.654717717717u,0 5803.655717717717u,1.5 5804.632257757758u,1.5 5804.633257757759u,0 5806.587337837837u,0 5806.588337837838u,1.5 5807.564877877878u,1.5 5807.565877877878u,0 5809.5199579579585u,0 5809.520957957959u,1.5 5811.475038038037u,1.5 5811.476038038038u,0 5812.452578078078u,0 5812.453578078078u,1.5 5814.4076581581585u,1.5 5814.408658158159u,0 5816.362738238237u,0 5816.363738238238u,1.5 5818.317818318318u,1.5 5818.318818318318u,0 5820.272898398398u,0 5820.273898398398u,1.5 5821.250438438438u,1.5 5821.2514384384385u,0 5822.227978478479u,0 5822.228978478479u,1.5 5827.115678678679u,1.5 5827.116678678679u,0 5834.935998998999u,0 5834.936998998999u,1.5 5836.891079079079u,1.5 5836.892079079079u,0 5837.868619119119u,0 5837.869619119119u,1.5 5839.823699199199u,1.5 5839.824699199199u,0 5842.756319319319u,0 5842.757319319319u,1.5 5843.7338593593595u,1.5 5843.73485935936u,0 5845.688939439439u,0 5845.6899394394395u,1.5 5846.66647947948u,1.5 5846.66747947948u,0 5847.644019519519u,0 5847.645019519519u,1.5 5849.5990995996u,1.5 5849.6000995996u,0 5850.576639639639u,0 5850.5776396396395u,1.5 5851.55417967968u,1.5 5851.55517967968u,0 5857.41941991992u,0 5857.42041991992u,1.5 5858.39695995996u,1.5 5858.397959959961u,0 5859.3745u,0 5859.3755u,1.5 5860.352040040039u,1.5 5860.35304004004u,0 5862.30712012012u,0 5862.30812012012u,1.5 5863.2846601601605u,1.5 5863.285660160161u,0 5864.2622002002u,0 5864.2632002002u,1.5 5865.239740240239u,1.5 5865.24074024024u,0 5866.217280280281u,0 5866.218280280281u,1.5 5867.19482032032u,1.5 5867.19582032032u,0 5871.104980480481u,0 5871.105980480481u,1.5 5872.08252052052u,1.5 5872.08352052052u,0 5873.0600605605605u,0 5873.061060560561u,1.5 5877.947760760761u,1.5 5877.948760760762u,0 5878.925300800801u,0 5878.926300800801u,1.5 5879.90284084084u,1.5 5879.9038408408405u,0 5880.880380880881u,0 5880.881380880881u,1.5 5881.857920920921u,1.5 5881.858920920921u,0 5882.835460960961u,0 5882.836460960962u,1.5 5883.813001001001u,1.5 5883.814001001001u,0 5885.768081081081u,0 5885.769081081081u,1.5 5888.700701201201u,1.5 5888.701701201201u,0 5889.67824124124u,0 5889.679241241241u,1.5 5891.633321321321u,1.5 5891.634321321321u,0 5892.6108613613615u,0 5892.611861361362u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5896.521021521521u,0 5896.522021521521u,1.5 5897.4985615615615u,1.5 5897.499561561562u,0 5899.453641641641u,0 5899.4546416416415u,1.5 5900.431181681682u,1.5 5900.432181681682u,0 5901.408721721721u,0 5901.409721721721u,1.5 5902.386261761762u,1.5 5902.387261761763u,0 5903.363801801802u,0 5903.364801801802u,1.5 5904.341341841841u,1.5 5904.3423418418415u,0 5905.318881881882u,0 5905.319881881882u,1.5 5907.273961961962u,1.5 5907.274961961963u,0 5908.251502002002u,0 5908.252502002002u,1.5 5910.206582082082u,1.5 5910.207582082082u,0 5911.184122122122u,0 5911.185122122122u,1.5 5913.139202202202u,1.5 5913.140202202202u,0 5921.9370625625625u,0 5921.938062562563u,1.5 5922.914602602603u,1.5 5922.915602602603u,0 5923.892142642642u,0 5923.8931426426425u,1.5 5926.824762762763u,1.5 5926.825762762764u,0 5927.802302802803u,0 5927.803302802803u,1.5 5930.734922922923u,1.5 5930.735922922923u,0 5931.712462962963u,0 5931.713462962964u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5942.465403403403u,0 5942.466403403403u,1.5 5944.420483483484u,1.5 5944.421483483484u,0 5945.398023523523u,0 5945.399023523523u,1.5 5946.375563563563u,1.5 5946.376563563564u,0 5949.308183683684u,0 5949.309183683684u,1.5 5950.285723723723u,1.5 5950.286723723723u,0 5952.240803803804u,0 5952.241803803804u,1.5 5953.218343843843u,1.5 5953.2193438438435u,0 5954.195883883884u,0 5954.196883883884u,1.5 5958.106044044043u,1.5 5958.1070440440435u,0 5959.083584084084u,0 5959.084584084084u,1.5 5962.993744244243u,1.5 5962.9947442442435u,0 5963.971284284285u,0 5963.972284284285u,1.5 5964.948824324324u,1.5 5964.949824324324u,0 5965.926364364364u,0 5965.927364364365u,1.5 5967.881444444444u,1.5 5967.882444444444u,0 5968.858984484485u,0 5968.859984484485u,1.5 5970.814064564564u,1.5 5970.815064564565u,0 5971.791604604605u,0 5971.792604604605u,1.5 5972.769144644644u,1.5 5972.7701446446445u,0 5973.746684684685u,0 5973.747684684685u,1.5 5974.724224724724u,1.5 5974.725224724724u,0 5976.679304804805u,0 5976.680304804805u,1.5 5977.656844844844u,1.5 5977.6578448448445u,0 5980.589464964965u,0 5980.590464964966u,1.5 5981.567005005005u,1.5 5981.568005005005u,0 5992.319945445445u,0 5992.320945445445u,1.5 5993.297485485486u,1.5 5993.298485485486u,0 5994.275025525525u,0 5994.276025525525u,1.5 5995.252565565565u,1.5 5995.253565565566u,0 5996.230105605606u,0 5996.231105605606u,1.5 5997.207645645645u,1.5 5997.208645645645u,0 6001.117805805806u,0 6001.118805805806u,1.5 6002.095345845845u,1.5 6002.0963458458455u,0 6013.825826326326u,0 6013.826826326326u,1.5 6014.803366366366u,1.5 6014.804366366367u,0 6019.691066566566u,0 6019.692066566567u,1.5 6020.668606606607u,1.5 6020.669606606607u,0 6024.578766766767u,0 6024.5797667667675u,1.5 6025.556306806807u,1.5 6025.557306806807u,0 6029.466466966967u,0 6029.467466966968u,1.5 6031.421547047046u,1.5 6031.4225470470465u,0 6035.331707207207u,0 6035.332707207207u,1.5 6036.309247247247u,1.5 6036.310247247247u,0 6038.264327327327u,0 6038.265327327327u,1.5 6045.107107607608u,1.5 6045.108107607608u,0 6046.084647647647u,0 6046.085647647647u,1.5 6048.039727727727u,1.5 6048.040727727727u,0 6049.017267767768u,0 6049.0182677677685u,1.5 6049.994807807808u,1.5 6049.995807807808u,0 6050.972347847847u,0 6050.973347847847u,1.5 6051.949887887888u,1.5 6051.950887887888u,0 6052.927427927928u,0 6052.928427927928u,1.5 6053.904967967968u,1.5 6053.9059679679685u,0 6061.7252882882885u,0 6061.726288288289u,1.5 6063.680368368368u,1.5 6063.681368368369u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6073.455768768769u,1.5 6073.4567687687695u,0 6077.365928928929u,0 6077.366928928929u,1.5 6078.343468968969u,1.5 6078.3444689689695u,0 6079.321009009009u,0 6079.322009009009u,1.5 6080.298549049048u,1.5 6080.299549049048u,0 6082.253629129129u,0 6082.254629129129u,1.5 6083.231169169169u,1.5 6083.2321691691695u,0 6084.208709209209u,0 6084.209709209209u,1.5 6085.186249249249u,1.5 6085.187249249249u,0 6087.141329329329u,0 6087.142329329329u,1.5 6088.118869369369u,1.5 6088.11986936937u,0 6090.073949449449u,0 6090.074949449449u,1.5 6091.0514894894895u,1.5 6091.05248948949u,0 6092.029029529529u,0 6092.030029529529u,1.5 6094.961649649649u,1.5 6094.962649649649u,0 6095.93918968969u,0 6095.94018968969u,1.5 6096.916729729729u,1.5 6096.917729729729u,0 6098.87180980981u,0 6098.87280980981u,1.5 6099.849349849849u,1.5 6099.850349849849u,0 6103.75951001001u,0 6103.76051001001u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6110.6022902902905u,1.5 6110.603290290291u,0 6111.57983033033u,0 6111.58083033033u,1.5 6114.51245045045u,1.5 6114.51345045045u,0 6116.46753053053u,0 6116.46853053053u,1.5 6117.44507057057u,1.5 6117.446070570571u,0 6120.3776906906905u,0 6120.378690690691u,1.5 6121.35523073073u,1.5 6121.35623073073u,0 6122.332770770771u,0 6122.3337707707715u,1.5 6123.310310810811u,1.5 6123.311310810811u,0 6124.28785085085u,0 6124.28885085085u,1.5 6128.198011011011u,1.5 6128.199011011011u,0 6129.17555105105u,0 6129.17655105105u,1.5 6130.1530910910915u,1.5 6130.154091091092u,0 6132.108171171171u,0 6132.1091711711715u,1.5 6134.063251251251u,1.5 6134.064251251251u,0 6136.995871371371u,0 6136.9968713713715u,1.5 6142.861111611612u,1.5 6142.862111611612u,0 6143.838651651651u,0 6143.839651651651u,1.5 6144.8161916916915u,1.5 6144.817191691692u,0 6147.748811811812u,0 6147.749811811812u,1.5 6148.726351851851u,1.5 6148.727351851851u,0 6149.7038918918915u,0 6149.704891891892u,1.5 6151.658971971972u,1.5 6151.6599719719725u,0 6152.636512012012u,0 6152.637512012012u,1.5 6156.546672172172u,1.5 6156.5476721721725u,0 6157.524212212212u,0 6157.525212212212u,1.5 6158.501752252252u,1.5 6158.502752252252u,0 6160.456832332332u,0 6160.457832332332u,1.5 6161.434372372372u,1.5 6161.4353723723725u,0 6162.411912412412u,0 6162.412912412412u,1.5 6163.389452452452u,1.5 6163.390452452452u,0 6164.3669924924925u,0 6164.367992492493u,1.5 6169.2546926926925u,1.5 6169.255692692693u,0 6170.232232732732u,0 6170.233232732732u,1.5 6171.209772772773u,1.5 6171.210772772773u,0 6172.187312812813u,0 6172.188312812813u,1.5 6173.164852852852u,1.5 6173.165852852852u,0 6175.119932932933u,0 6175.120932932933u,1.5 6180.985173173173u,1.5 6180.9861731731735u,0 6186.850413413413u,0 6186.851413413413u,1.5 6190.760573573573u,1.5 6190.7615735735735u,0 6195.648273773774u,0 6195.649273773774u,1.5 6196.625813813814u,1.5 6196.626813813814u,0 6197.603353853853u,0 6197.604353853853u,1.5 6202.491054054053u,1.5 6202.492054054053u,0 6207.378754254254u,0 6207.379754254254u,1.5 6213.2439944944945u,1.5 6213.244994494495u,0 6214.221534534534u,0 6214.222534534534u,1.5 6215.199074574574u,1.5 6215.2000745745745u,0 6217.154154654654u,0 6217.155154654654u,1.5 6219.109234734734u,1.5 6219.110234734734u,0 6220.086774774775u,0 6220.087774774775u,1.5 6223.0193948948945u,1.5 6223.020394894895u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6230.839715215215u,1.5 6230.840715215215u,0 6231.817255255255u,0 6231.818255255255u,1.5 6234.749875375375u,1.5 6234.7508753753755u,0 6238.660035535535u,0 6238.661035535535u,1.5 6239.637575575575u,1.5 6239.6385755755755u,0 6240.615115615616u,0 6240.616115615616u,1.5 6244.525275775776u,1.5 6244.526275775776u,0 6247.4578958958955u,0 6247.458895895896u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6252.345596096096u,0 6252.346596096097u,1.5 6253.323136136136u,1.5 6253.324136136136u,0 6255.278216216216u,0 6255.279216216216u,1.5 6256.255756256256u,1.5 6256.256756256256u,0 6257.233296296296u,0 6257.234296296297u,1.5 6258.210836336336u,1.5 6258.211836336336u,0 6259.188376376376u,0 6259.1893763763765u,1.5 6260.165916416417u,1.5 6260.166916416417u,0 6261.143456456457u,0 6261.144456456457u,1.5 6262.120996496496u,1.5 6262.121996496497u,0 6263.098536536536u,0 6263.099536536536u,1.5 6268.963776776777u,1.5 6268.964776776777u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6274.829017017017u,1.5 6274.830017017017u,0 6275.806557057057u,0 6275.807557057057u,1.5 6276.784097097097u,1.5 6276.785097097098u,0 6277.761637137137u,0 6277.762637137137u,1.5 6278.739177177177u,1.5 6278.740177177177u,0 6279.716717217217u,0 6279.717717217217u,1.5 6280.694257257258u,1.5 6280.695257257258u,0 6281.671797297297u,0 6281.672797297298u,1.5 6282.649337337337u,1.5 6282.650337337337u,0 6283.626877377377u,0 6283.627877377377u,1.5 6285.581957457458u,1.5 6285.582957457458u,0 6286.559497497497u,0 6286.560497497498u,1.5 6287.537037537537u,1.5 6287.538037537537u,0 6288.514577577577u,0 6288.5155775775775u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6293.402277777778u,0 6293.403277777778u,1.5 6296.3348978978975u,1.5 6296.335897897898u,0 6297.312437937938u,0 6297.313437937938u,1.5 6299.267518018018u,1.5 6299.268518018018u,0 6300.245058058058u,0 6300.246058058058u,1.5 6301.222598098098u,1.5 6301.223598098099u,0 6303.177678178178u,0 6303.178678178178u,1.5 6307.087838338338u,1.5 6307.088838338338u,0 6308.065378378378u,0 6308.066378378378u,1.5 6309.042918418419u,1.5 6309.043918418419u,0 6310.997998498498u,0 6310.998998498499u,1.5 6311.975538538538u,1.5 6311.976538538538u,0 6315.885698698698u,0 6315.886698698699u,1.5 6320.773398898898u,1.5 6320.774398898899u,0 6322.728478978979u,0 6322.729478978979u,1.5 6324.683559059059u,1.5 6324.684559059059u,0 6325.661099099099u,0 6325.6620990991u,1.5 6326.638639139139u,1.5 6326.639639139139u,0 6327.616179179179u,0 6327.617179179179u,1.5 6330.548799299299u,1.5 6330.5497992993u,0 6331.526339339339u,0 6331.527339339339u,1.5 6332.503879379379u,1.5 6332.504879379379u,0 6338.36911961962u,0 6338.37011961962u,1.5 6344.23435985986u,1.5 6344.23535985986u,0 6345.211899899899u,0 6345.2128998999u,1.5 6346.18943993994u,1.5 6346.19043993994u,0 6347.16697997998u,0 6347.16797997998u,1.5 6348.14452002002u,1.5 6348.14552002002u,0 6350.0996001001u,0 6350.100600100101u,1.5 6351.07714014014u,1.5 6351.07814014014u,0 6352.05468018018u,0 6352.05568018018u,1.5 6355.96484034034u,1.5 6355.96584034034u,0 6359.8750005005u,0 6359.876000500501u,1.5 6360.85254054054u,1.5 6360.85354054054u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6364.7627007007u,0 6364.763700700701u,1.5 6367.695320820821u,1.5 6367.696320820821u,0 6369.6504009009u,0 6369.651400900901u,1.5 6370.627940940941u,1.5 6370.628940940941u,0 6372.583021021021u,0 6372.584021021021u,1.5 6373.560561061061u,1.5 6373.561561061061u,0 6374.538101101101u,0 6374.539101101102u,1.5 6376.493181181181u,1.5 6376.494181181181u,0 6378.448261261262u,0 6378.449261261262u,1.5 6381.380881381381u,1.5 6381.381881381381u,0 6383.335961461462u,0 6383.336961461462u,1.5 6386.268581581581u,1.5 6386.269581581581u,0 6389.201201701701u,0 6389.202201701702u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6393.111361861862u,0 6393.112361861862u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6396.043981981982u,1.5 6396.044981981982u,0 6397.021522022022u,0 6397.022522022022u,1.5 6399.954142142142u,1.5 6399.955142142142u,0 6400.931682182182u,0 6400.932682182182u,1.5 6402.886762262263u,1.5 6402.887762262263u,0 6403.864302302302u,0 6403.865302302303u,1.5 6404.841842342342u,1.5 6404.842842342342u,0 6411.684622622623u,0 6411.685622622623u,1.5 6412.662162662663u,1.5 6412.663162662663u,0 6413.639702702702u,0 6413.640702702703u,1.5 6414.617242742742u,1.5 6414.618242742742u,0 6416.572322822823u,0 6416.573322822823u,1.5 6419.504942942943u,1.5 6419.505942942943u,0 6421.460023023023u,0 6421.461023023023u,1.5 6422.437563063063u,1.5 6422.438563063063u,0 6427.325263263264u,0 6427.326263263264u,1.5 6428.302803303303u,1.5 6428.3038033033035u,0 6432.212963463464u,0 6432.213963463464u,1.5 6433.190503503503u,1.5 6433.191503503504u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6436.1231236236235u,0 6436.124123623624u,1.5 6438.078203703703u,1.5 6438.079203703704u,0 6439.055743743743u,0 6439.056743743743u,1.5 6442.965903903903u,1.5 6442.966903903904u,0 6443.943443943944u,0 6443.944443943944u,1.5 6446.876064064064u,1.5 6446.877064064064u,0 6447.853604104104u,0 6447.8546041041045u,1.5 6448.831144144144u,1.5 6448.832144144144u,0 6449.808684184184u,0 6449.809684184184u,1.5 6450.786224224224u,1.5 6450.787224224224u,0 6451.763764264265u,0 6451.764764264265u,1.5 6452.741304304304u,1.5 6452.7423043043045u,0 6456.651464464465u,0 6456.652464464465u,1.5 6457.629004504504u,1.5 6457.6300045045045u,0 6460.5616246246245u,0 6460.562624624625u,1.5 6461.539164664665u,1.5 6461.540164664665u,0 6466.426864864865u,0 6466.427864864865u,1.5 6467.404404904904u,1.5 6467.405404904905u,0 6468.381944944945u,0 6468.382944944945u,1.5 6469.359484984985u,1.5 6469.360484984985u,0 6470.337025025025u,0 6470.338025025025u,1.5 6471.314565065065u,1.5 6471.315565065065u,0 6472.292105105105u,0 6472.2931051051055u,1.5 6473.269645145145u,1.5 6473.270645145145u,0 6474.247185185185u,0 6474.248185185185u,1.5 6477.179805305305u,1.5 6477.1808053053055u,0 6478.157345345345u,0 6478.158345345345u,1.5 6483.045045545545u,1.5 6483.046045545545u,0 6485.977665665666u,0 6485.978665665666u,1.5 6486.955205705705u,1.5 6486.9562057057055u,0 6487.932745745745u,0 6487.933745745745u,1.5 6489.8878258258255u,1.5 6489.888825825826u,0 6491.842905905905u,0 6491.843905905906u,1.5 6494.775526026026u,1.5 6494.776526026026u,0 6496.730606106106u,0 6496.7316061061065u,1.5 6500.640766266267u,1.5 6500.641766266267u,0 6501.618306306306u,0 6501.6193063063065u,1.5 6502.595846346346u,1.5 6502.596846346346u,0 6505.528466466467u,0 6505.529466466467u,1.5 6508.461086586587u,1.5 6508.462086586587u,0 6510.416166666667u,0 6510.417166666667u,1.5 6512.371246746747u,1.5 6512.372246746747u,0 6515.303866866867u,0 6515.304866866867u,1.5 6516.281406906906u,1.5 6516.2824069069065u,0 6517.258946946947u,0 6517.259946946947u,1.5 6519.2140270270265u,1.5 6519.215027027027u,0 6520.191567067067u,0 6520.192567067067u,1.5 6521.169107107107u,1.5 6521.1701071071075u,0 6522.146647147147u,0 6522.147647147147u,1.5 6523.124187187187u,1.5 6523.125187187187u,0 6524.101727227227u,0 6524.102727227227u,1.5 6525.079267267268u,1.5 6525.080267267268u,0 6526.056807307307u,0 6526.0578073073075u,1.5 6528.011887387387u,1.5 6528.012887387387u,0 6529.966967467468u,0 6529.967967467468u,1.5 6531.922047547547u,1.5 6531.923047547547u,0 6532.899587587588u,0 6532.900587587588u,1.5 6533.8771276276275u,1.5 6533.878127627628u,0 6534.854667667668u,0 6534.855667667668u,1.5 6535.832207707707u,1.5 6535.8332077077075u,0 6536.809747747748u,0 6536.810747747748u,1.5 6537.787287787788u,1.5 6537.788287787788u,0 6538.7648278278275u,0 6538.765827827828u,1.5 6539.742367867868u,1.5 6539.743367867868u,0 6545.607608108108u,0 6545.6086081081085u,1.5 6546.585148148148u,1.5 6546.586148148148u,0 6547.562688188188u,0 6547.563688188188u,1.5 6548.5402282282275u,1.5 6548.541228228228u,0 6550.495308308308u,0 6550.4963083083085u,1.5 6552.450388388388u,1.5 6552.451388388388u,0 6553.4279284284285u,0 6553.428928428429u,1.5 6554.405468468469u,1.5 6554.406468468469u,0 6555.383008508508u,0 6555.3840085085085u,1.5 6556.360548548548u,1.5 6556.361548548548u,0 6558.3156286286285u,0 6558.316628628629u,1.5 6560.270708708708u,1.5 6560.2717087087085u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6566.135948948949u,0 6566.136948948949u,1.5 6567.113488988989u,1.5 6567.114488988989u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.9787292292285u,1.5 6572.979729229229u,0 6573.95626926927u,0 6573.95726926927u,1.5 6575.911349349349u,1.5 6575.912349349349u,0 6577.866429429429u,0 6577.86742942943u,1.5 6578.84396946947u,1.5 6578.84496946947u,0 6579.821509509509u,0 6579.8225095095095u,1.5 6584.709209709709u,1.5 6584.7102097097095u,0 6588.61936986987u,0 6588.62036986987u,1.5 6592.5295300300295u,1.5 6592.53053003003u,0 6598.394770270271u,0 6598.395770270271u,1.5 6599.37231031031u,1.5 6599.37331031031u,0 6601.32739039039u,0 6601.32839039039u,1.5 6602.30493043043u,1.5 6602.305930430431u,0 6603.282470470471u,0 6603.283470470471u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6608.170170670671u,0 6608.171170670671u,1.5 6609.14771071071u,1.5 6609.1487107107105u,0 6614.03541091091u,0 6614.0364109109105u,1.5 6615.990490990991u,1.5 6615.991490990991u,0 6616.9680310310305u,0 6616.969031031031u,1.5 6619.900651151151u,1.5 6619.901651151151u,0 6620.878191191191u,0 6620.879191191191u,1.5 6622.833271271272u,1.5 6622.834271271272u,0 6623.810811311311u,0 6623.811811311311u,1.5 6624.788351351351u,1.5 6624.789351351351u,0 6629.676051551551u,0 6629.677051551551u,1.5 6630.653591591592u,1.5 6630.654591591592u,0 6633.586211711711u,0 6633.5872117117115u,1.5 6634.563751751752u,1.5 6634.564751751752u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6640.428991991992u,0 6640.429991991992u,1.5 6642.384072072072u,1.5 6642.385072072072u,0 6643.361612112112u,0 6643.362612112112u,1.5 6645.316692192192u,1.5 6645.317692192192u,0 6646.2942322322315u,0 6646.295232232232u,1.5 6650.204392392392u,1.5 6650.205392392392u,0 6652.159472472473u,0 6652.160472472473u,1.5 6654.114552552552u,1.5 6654.115552552552u,0 6655.092092592593u,0 6655.093092592593u,1.5 6656.069632632632u,1.5 6656.070632632633u,0 6657.047172672673u,0 6657.048172672673u,1.5 6658.024712712712u,1.5 6658.025712712712u,0 6659.002252752753u,0 6659.003252752753u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6666.822573073073u,0 6666.823573073073u,1.5 6667.800113113113u,1.5 6667.801113113113u,0 6668.777653153153u,0 6668.778653153153u,1.5 6671.710273273274u,1.5 6671.711273273274u,0 6672.687813313313u,0 6672.688813313313u,1.5 6674.642893393393u,1.5 6674.643893393393u,0 6676.597973473474u,0 6676.598973473474u,1.5 6677.575513513513u,1.5 6677.576513513513u,0 6678.553053553553u,0 6678.554053553553u,1.5 6679.530593593594u,1.5 6679.531593593594u,0 6680.508133633633u,0 6680.509133633634u,1.5 6684.418293793794u,1.5 6684.419293793794u,0 6685.395833833833u,0 6685.396833833834u,1.5 6687.350913913913u,1.5 6687.351913913913u,0 6689.305993993994u,0 6689.306993993994u,1.5 6690.283534034033u,1.5 6690.284534034034u,0 6692.238614114114u,0 6692.239614114114u,1.5 6697.126314314314u,1.5 6697.127314314314u,0 6702.991554554554u,0 6702.992554554554u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6710.811874874875u,0 6710.812874874875u,1.5 6711.789414914914u,1.5 6711.790414914914u,0 6712.766954954955u,0 6712.767954954955u,1.5 6713.744494994995u,1.5 6713.745494994995u,0 6714.722035035034u,0 6714.723035035035u,1.5 6715.699575075075u,1.5 6715.700575075075u,0 6717.654655155155u,0 6717.655655155155u,1.5 6719.609735235234u,1.5 6719.610735235235u,0 6720.587275275276u,0 6720.588275275276u,1.5 6724.497435435435u,1.5 6724.498435435436u,0 6726.452515515515u,0 6726.453515515515u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6730.362675675676u,0 6730.363675675676u,1.5 6731.340215715715u,1.5 6731.341215715715u,0 6734.272835835835u,0 6734.273835835836u,1.5 6735.250375875876u,1.5 6735.251375875876u,0 6736.227915915916u,0 6736.228915915916u,1.5 6739.160536036035u,1.5 6739.161536036036u,0 6740.138076076076u,0 6740.139076076076u,1.5 6741.115616116116u,1.5 6741.116616116116u,0 6742.093156156156u,0 6742.094156156156u,1.5 6743.070696196196u,1.5 6743.071696196196u,0 6745.025776276277u,0 6745.026776276277u,1.5 6746.980856356356u,1.5 6746.981856356356u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6755.778716716716u,0 6755.779716716716u,1.5 6756.7562567567575u,1.5 6756.757256756758u,0 6759.688876876877u,0 6759.689876876877u,1.5 6762.621496996997u,1.5 6762.622496996997u,0 6766.5316571571575u,0 6766.532657157158u,1.5 6770.441817317317u,1.5 6770.442817317317u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6776.3070575575575u,0 6776.308057557558u,1.5 6780.217217717717u,1.5 6780.218217717717u,0 6784.127377877878u,0 6784.128377877878u,1.5 6785.104917917918u,1.5 6785.105917917918u,0 6788.037538038037u,0 6788.038538038038u,1.5 6792.925238238237u,1.5 6792.926238238238u,0 6798.790478478479u,0 6798.791478478479u,1.5 6799.768018518518u,1.5 6799.769018518518u,0 6800.7455585585585u,0 6800.746558558559u,1.5 6802.700638638638u,1.5 6802.7016386386385u,0 6804.655718718718u,0 6804.656718718718u,1.5 6806.610798798799u,1.5 6806.611798798799u,0 6808.565878878879u,0 6808.566878878879u,1.5 6809.543418918919u,1.5 6809.544418918919u,0 6810.520958958959u,0 6810.52195895896u,1.5 6812.476039039038u,1.5 6812.477039039039u,0 6813.453579079079u,0 6813.454579079079u,1.5 6816.386199199199u,1.5 6816.387199199199u,0 6819.318819319319u,0 6819.319819319319u,1.5 6820.2963593593595u,1.5 6820.29735935936u,0 6821.273899399399u,0 6821.274899399399u,1.5 6823.22897947948u,1.5 6823.22997947948u,0 6825.1840595595595u,0 6825.18505955956u,1.5 6826.1615995996u,1.5 6826.1625995996u,0 6827.139139639639u,0 6827.1401396396395u,1.5 6828.11667967968u,1.5 6828.11767967968u,0 6831.0492997998u,0 6831.0502997998u,1.5 6832.026839839839u,1.5 6832.0278398398395u,0 6833.00437987988u,0 6833.00537987988u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6843.75732032032u,0 6843.75832032032u,1.5 6844.7348603603605u,1.5 6844.735860360361u,0 6845.7124004004u,0 6845.7134004004u,1.5 6846.68994044044u,1.5 6846.6909404404405u,0 6847.667480480481u,0 6847.668480480481u,1.5 6850.600100600601u,1.5 6850.601100600601u,0 6854.510260760761u,0 6854.511260760762u,1.5 6855.487800800801u,1.5 6855.488800800801u,0 6856.46534084084u,0 6856.4663408408405u,1.5 6857.442880880881u,1.5 6857.443880880881u,0 6859.397960960961u,0 6859.398960960962u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6865.263201201201u,0 6865.264201201201u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6872.105981481482u,0 6872.106981481482u,1.5 6873.083521521521u,1.5 6873.084521521521u,0 6874.0610615615615u,0 6874.062061561562u,1.5 6877.971221721721u,1.5 6877.972221721721u,0 6878.948761761762u,0 6878.949761761763u,1.5 6879.926301801802u,1.5 6879.927301801802u,0 6883.836461961962u,0 6883.837461961963u,1.5 6884.814002002002u,1.5 6884.815002002002u,0 6886.769082082082u,0 6886.770082082082u,1.5 6889.701702202202u,1.5 6889.702702202202u,0 6890.679242242241u,0 6890.680242242242u,1.5 6891.656782282283u,1.5 6891.657782282283u,0 6892.634322322322u,0 6892.635322322322u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6902.409722722722u,0 6902.410722722722u,1.5 6903.387262762763u,1.5 6903.388262762764u,0 6904.364802802803u,0 6904.365802802803u,1.5 6911.207583083083u,1.5 6911.208583083083u,0 6912.185123123123u,0 6912.186123123123u,1.5 6913.162663163163u,1.5 6913.163663163164u,0 6915.117743243242u,0 6915.1187432432425u,1.5 6916.095283283284u,1.5 6916.096283283284u,0 6918.050363363363u,0 6918.051363363364u,1.5 6919.027903403403u,1.5 6919.028903403403u,0 6921.960523523523u,0 6921.961523523523u,1.5 6924.893143643643u,1.5 6924.8941436436435u,0 6925.870683683684u,0 6925.871683683684u,1.5 6929.780843843843u,1.5 6929.7818438438435u,0 6930.758383883884u,0 6930.759383883884u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6937.601164164164u,0 6937.602164164165u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6943.466404404404u,0 6943.467404404404u,1.5 6945.421484484485u,1.5 6945.422484484485u,0 6946.399024524524u,0 6946.400024524524u,1.5 6947.376564564564u,1.5 6947.377564564565u,0 6949.331644644644u,0 6949.3326446446445u,1.5 6952.264264764765u,1.5 6952.265264764766u,0 6953.241804804805u,0 6953.242804804805u,1.5 6956.174424924925u,1.5 6956.175424924925u,0 6959.107045045044u,0 6959.1080450450445u,1.5 6963.994745245244u,1.5 6963.9957452452445u,0 6964.972285285286u,0 6964.973285285286u,1.5 6965.949825325325u,1.5 6965.950825325325u,0 6966.927365365365u,0 6966.928365365366u,1.5 6968.882445445445u,1.5 6968.883445445445u,0 6971.815065565565u,0 6971.816065565566u,1.5 6972.792605605606u,1.5 6972.793605605606u,0 6973.770145645645u,0 6973.771145645645u,1.5 6974.747685685686u,1.5 6974.748685685686u,0 6975.725225725725u,0 6975.726225725725u,1.5 6976.702765765766u,1.5 6976.703765765767u,0 6980.612925925926u,0 6980.613925925926u,1.5 6981.590465965966u,1.5 6981.591465965967u,0 6986.478166166166u,0 6986.479166166167u,1.5 6989.410786286287u,1.5 6989.411786286287u,0 6990.388326326326u,0 6990.389326326326u,1.5 6991.365866366366u,1.5 6991.366866366367u,0 6992.343406406406u,0 6992.344406406406u,1.5 6993.320946446446u,1.5 6993.321946446446u,0 6996.253566566566u,0 6996.254566566567u,1.5 6997.231106606607u,1.5 6997.232106606607u,0
vbb22 bb22 0 pwl 0,1.5  17.59522072072072u,1.5 17.59622072072072u,0 18.572760760760765u,0 18.573760760760763u,1.5 21.50538088088088u,1.5 21.50638088088088u,0 22.482920920920925u,0 22.483920920920923u,1.5 27.370621121121122u,1.5 27.37162112112112u,0 28.348161161161162u,0 28.34916116116116u,1.5 29.325701201201202u,1.5 29.3267012012012u,0 30.303241241241246u,0 30.304241241241243u,1.5 32.25832132132132u,1.5 32.25932132132132u,0 37.146021521521526u,0 37.14702152152153u,1.5 38.12356156156156u,1.5 38.12456156156156u,0 40.07864164164164u,0 40.07964164164164u,1.5 41.05618168168168u,1.5 41.05718168168168u,0 61.58452252252251u,0 61.58552252252252u,1.5 62.56206256256256u,1.5 62.563062562562564u,0 63.539602602602606u,0 63.54060260260261u,1.5 64.51714264264264u,1.5 64.51814264264264u,0 65.49468268268268u,0 65.49568268268268u,1.5 66.47222272272272u,1.5 66.47322272272272u,0 67.44976276276276u,0 67.45076276276276u,1.5 68.4273028028028u,1.5 68.4283028028028u,0 69.40484284284284u,0 69.40584284284284u,1.5 70.38238288288288u,1.5 70.38338288288288u,0 71.35992292292292u,0 71.36092292292292u,1.5 81.13532332332332u,1.5 81.13632332332332u,0 82.11286336336336u,0 82.11386336336336u,1.5 85.04548348348348u,1.5 85.04648348348348u,0 86.02302352352352u,0 86.02402352352352u,1.5 88.95564364364364u,1.5 88.95664364364364u,0 89.9331836836837u,0 89.9341836836837u,1.5 90.91072372372372u,1.5 90.91172372372372u,0 107.5289044044044u,0 107.5299044044044u,1.5 120.23692492492492u,1.5 120.23792492492493u,0 121.21446496496498u,0 121.21546496496498u,1.5 122.19200500500502u,1.5 122.19300500500502u,0 124.14708508508508u,0 124.14808508508509u,1.5 125.12462512512512u,1.5 125.12562512512513u,0 134.90002552552554u,0 134.9010255255255u,1.5 135.8775655655656u,1.5 135.87856556556557u,0 137.83264564564567u,0 137.83364564564565u,1.5 148.58558608608612u,1.5 148.5865860860861u,0 149.56312612612612u,0 149.5641261261261u,1.5 150.54066616616618u,1.5 150.54166616616615u,0 151.51820620620623u,0 151.5192062062062u,1.5 152.49574624624626u,1.5 152.49674624624623u,0 163.2486866866867u,0 163.2496866866867u,1.5 174.00162712712714u,1.5 174.0026271271271u,0 177.9117872872873u,0 177.91278728728727u,1.5 178.88932732732735u,1.5 178.89032732732733u,0 184.7545675675676u,0 184.75556756756757u,1.5 186.70964764764764u,1.5 186.71064764764762u,0 187.6871876876877u,0 187.68818768768767u,1.5 194.529967967968u,1.5 194.53096796796797u,0 195.50750800800802u,0 195.508508008008u,1.5 197.4625880880881u,1.5 197.46358808808807u,0 208.21552852852852u,0 208.2165285285285u,1.5 217.0133888888889u,1.5 217.01438888888887u,0 217.99092892892892u,0 217.9919289289289u,1.5 218.96846896896898u,1.5 218.96946896896895u,0 221.90108908908908u,0 221.90208908908906u,1.5 222.87862912912914u,1.5 222.8796291291291u,0 225.81124924924927u,0 225.81224924924925u,1.5 226.7887892892893u,1.5 226.78978928928927u,0 228.74386936936938u,0 228.74486936936935u,1.5 239.4968098098098u,1.5 239.49780980980978u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 259.04761061061066u,1.5 259.04861061061064u,0 260.02515065065063u,0 260.0261506506506u,1.5 261.98023073073074u,1.5 261.9812307307307u,0 262.95777077077076u,0 262.95877077077074u,1.5 263.93531081081085u,1.5 263.9363108108108u,0 264.9128508508509u,0 264.91385085085085u,1.5 265.8903908908909u,1.5 265.8913908908909u,0 271.75563113113117u,0 271.75663113113114u,1.5 280.5534914914915u,1.5 280.5544914914915u,0 281.53103153153154u,0 281.5320315315315u,1.5 282.50857157157157u,1.5 282.50957157157154u,0 283.48611161161165u,0 283.4871116116116u,1.5 284.4636516516517u,1.5 284.46465165165165u,0 291.3064319319319u,0 291.3074319319319u,1.5 292.28397197197194u,1.5 292.2849719719719u,0 294.23905205205205u,0 294.240052052052u,1.5 302.0593723723724u,1.5 302.0603723723724u,0 303.03691241241245u,0 303.0379124124124u,1.5 304.9919924924925u,1.5 304.9929924924925u,0 314.76739289289293u,0 314.7683928928929u,1.5 316.722472972973u,1.5 316.72347297297296u,0 317.700013013013u,0 317.701013013013u,1.5 325.5203333333333u,1.5 325.5213333333333u,0 326.4978733733734u,0 326.4988733733734u,1.5 327.47541341341343u,1.5 327.4764134134134u,0 329.4304934934935u,0 329.43149349349346u,1.5 330.4080335335335u,1.5 330.4090335335335u,0 334.31819369369373u,0 334.3191936936937u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 337.2508138138138u,0 337.2518138138138u,1.5 348.9812942942943u,1.5 348.98229429429426u,0 349.9588343343343u,0 349.9598343343343u,1.5 350.9363743743744u,1.5 350.9373743743744u,0 351.9139144144144u,0 351.9149144144144u,1.5 352.8914544544545u,1.5 352.8924544544545u,0 353.8689944944945u,0 353.86999449449445u,1.5 354.8465345345345u,1.5 354.8475345345345u,0 362.6668548548549u,0 362.66785485485485u,1.5 363.6443948948949u,1.5 363.6453948948949u,0 364.621934934935u,0 364.62293493493496u,1.5 377.3299554554555u,1.5 377.33095545545547u,0 378.3074954954955u,0 378.3084954954955u,1.5 379.28503553553554u,1.5 379.2860355355355u,0 391.99305605605605u,0 391.994056056056u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 406.65615665665666u,1.5 406.65715665665664u,0 407.6336966966967u,0 407.63469669669666u,1.5 409.5887767767768u,1.5 409.5897767767768u,0 410.5663168168168u,0 410.5673168168168u,1.5 413.49893693693696u,1.5 413.49993693693693u,0 416.43155705705703u,0 416.432557057057u,1.5 417.40909709709706u,1.5 417.41009709709704u,0 434.0272777777778u,0 434.02827777777776u,1.5 435.98235785785783u,1.5 435.9833578578578u,0 436.9598978978979u,0 436.9608978978979u,1.5 442.82513813813813u,1.5 442.8261381381381u,0 443.80267817817816u,0 443.80367817817813u,1.5 447.7128383383383u,1.5 447.7138383383383u,0 448.69037837837834u,0 448.6913783783783u,1.5 462.37593893893893u,1.5 462.3769389389389u,0 463.353478978979u,0 463.354478978979u,1.5 467.2636391391391u,1.5 467.2646391391391u,0 468.2411791791792u,0 468.2421791791792u,1.5 470.19625925925925u,1.5 470.1972592592592u,0 472.15133933933936u,0 472.15233933933933u,1.5 473.1288793793794u,1.5 473.12987937937936u,0 474.1064194194194u,0 474.1074194194194u,1.5 475.08395945945944u,1.5 475.0849594594594u,0 478.0165795795796u,0 478.0175795795796u,1.5 478.9941196196196u,1.5 478.9951196196196u,0 481.92673973973973u,0 481.9277397397397u,1.5 482.9042797797798u,1.5 482.9052797797798u,0 484.8593598598599u,0 484.8603598598599u,1.5 485.8368998998999u,1.5 485.83789989989987u,0 489.7470600600601u,0 489.7480600600601u,1.5 490.72460010010013u,1.5 490.7256001001001u,0 512.2304809809809u,0 512.2314809809809u,1.5 513.2080210210211u,1.5 513.209021021021u,0 514.1855610610611u,0 514.1865610610611u,1.5 515.1631011011011u,1.5 515.1641011011011u,0 516.1406411411411u,0 516.1416411411411u,1.5 517.1181811811812u,1.5 517.1191811811811u,0 518.0957212212213u,0 518.0967212212213u,1.5 519.0732612612613u,1.5 519.0742612612613u,0 520.0508013013012u,0 520.0518013013012u,1.5 521.0283413413413u,1.5 521.0293413413413u,0 525.9160415415415u,0 525.9170415415415u,1.5 526.8935815815815u,1.5 526.8945815815815u,0 527.8711216216217u,0 527.8721216216217u,1.5 529.8262017017017u,1.5 529.8272017017017u,0 531.7812817817818u,0 531.7822817817818u,1.5 534.7139019019019u,1.5 534.7149019019018u,0 535.6914419419419u,0 535.6924419419419u,1.5 537.646522022022u,1.5 537.647522022022u,0 538.6240620620621u,0 538.625062062062u,1.5 560.1299429429429u,1.5 560.1309429429429u,0 562.085023023023u,0 562.086023023023u,1.5 565.0176431431431u,1.5 565.0186431431431u,0 565.9951831831833u,0 565.9961831831832u,1.5 566.9727232232233u,1.5 566.9737232232233u,0 567.9502632632633u,0 567.9512632632633u,1.5 568.9278033033033u,1.5 568.9288033033033u,0 587.501064064064u,0 587.502064064064u,1.5 588.4786041041041u,1.5 588.479604104104u,0 589.4561441441441u,0 589.4571441441441u,1.5 591.4112242242243u,1.5 591.4122242242242u,0 592.3887642642643u,0 592.3897642642643u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 607.0518648648649u,0 607.0528648648649u,1.5 608.0294049049048u,1.5 608.0304049049048u,0 619.7598853853854u,0 619.7608853853853u,1.5 620.7374254254254u,1.5 620.7384254254254u,0 621.7149654654654u,0 621.7159654654654u,1.5 622.6925055055054u,1.5 622.6935055055054u,0 623.6700455455456u,0 623.6710455455456u,1.5 633.445445945946u,1.5 633.4464459459459u,0 634.422985985986u,0 634.423985985986u,1.5 635.400526026026u,1.5 635.401526026026u,0 636.378066066066u,0 636.379066066066u,1.5 637.355606106106u,1.5 637.356606106106u,0 646.1534664664664u,0 646.1544664664664u,1.5 647.1310065065064u,1.5 647.1320065065064u,0 650.0636266266266u,0 650.0646266266266u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 664.7267272272272u,0 664.7277272272272u,1.5 665.7042672672673u,1.5 665.7052672672672u,0 673.5245875875876u,0 673.5255875875876u,1.5 674.5021276276276u,1.5 674.5031276276276u,0 675.4796676676676u,0 675.4806676676676u,1.5 678.4122877877878u,1.5 678.4132877877878u,0 679.3898278278278u,0 679.3908278278278u,1.5 684.277528028028u,1.5 684.278528028028u,0 687.2101481481482u,0 687.2111481481481u,1.5 688.1876881881882u,1.5 688.1886881881882u,0 696.9855485485485u,0 696.9865485485485u,1.5 697.9630885885886u,1.5 697.9640885885885u,0 698.9406286286286u,0 698.9416286286286u,1.5 704.8058688688689u,1.5 704.8068688688688u,0 705.783408908909u,0 705.784408908909u,1.5 708.716029029029u,1.5 708.7170290290289u,0 718.4914294294294u,0 718.4924294294294u,1.5 719.4689694694696u,1.5 719.4699694694696u,0 720.4465095095095u,0 720.4475095095095u,1.5 727.2892897897898u,1.5 727.2902897897898u,0 728.2668298298298u,0 728.2678298298298u,1.5 730.22190990991u,1.5 730.22290990991u,0 739.0197702702703u,0 739.0207702702703u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 758.5705710710711u,0 758.571571071071u,1.5 759.5481111111111u,1.5 759.5491111111111u,0 761.5031911911911u,0 761.5041911911911u,1.5 763.4582712712713u,1.5 763.4592712712713u,0 764.4358113113113u,0 764.4368113113113u,1.5 770.3010515515515u,1.5 770.3020515515515u,0 780.076451951952u,0 780.077451951952u,1.5 781.053991991992u,1.5 781.054991991992u,0 783.0090720720721u,0 783.010072072072u,1.5 791.8069324324325u,1.5 791.8079324324325u,0 801.5823328328329u,0 801.5833328328329u,1.5 802.5598728728729u,1.5 802.5608728728729u,0 803.5374129129129u,0 803.5384129129129u,1.5 804.514952952953u,1.5 804.515952952953u,0 805.492492992993u,0 805.493492992993u,1.5 813.3128133133133u,1.5 813.3138133133133u,0 815.2678933933934u,0 815.2688933933933u,1.5 816.2454334334335u,1.5 816.2464334334335u,0 817.2229734734735u,0 817.2239734734735u,1.5 818.2005135135136u,1.5 818.2015135135135u,0 825.0432937937937u,0 825.0442937937937u,1.5 826.0208338338339u,1.5 826.0218338338339u,0 826.9983738738739u,0 826.9993738738739u,1.5 834.8186941941941u,1.5 834.8196941941941u,0 835.7962342342342u,0 835.7972342342342u,1.5 836.7737742742743u,1.5 836.7747742742743u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 849.4817947947948u,0 849.4827947947948u,1.5 850.4593348348349u,1.5 850.4603348348348u,0 851.4368748748749u,0 851.4378748748749u,1.5 853.3919549549549u,1.5 853.3929549549549u,0 854.3694949949951u,0 854.370494994995u,1.5 861.2122752752753u,1.5 861.2132752752752u,0 862.1898153153153u,0 862.1908153153153u,1.5 863.1673553553553u,1.5 863.1683553553553u,0 865.1224354354355u,0 865.1234354354355u,1.5 866.0999754754755u,1.5 866.1009754754755u,0 874.8978358358358u,0 874.8988358358358u,1.5 875.8753758758759u,1.5 875.8763758758759u,0 877.8304559559559u,0 877.8314559559559u,1.5 878.8079959959961u,1.5 878.808995995996u,0 879.7855360360361u,0 879.7865360360361u,1.5 895.4261766766766u,1.5 895.4271766766766u,0 905.2015770770771u,0 905.2025770770771u,1.5 906.1791171171171u,1.5 906.1801171171171u,0 910.0892772772772u,0 910.0902772772772u,1.5 911.0668173173173u,1.5 911.0678173173172u,0 912.0443573573574u,0 912.0453573573574u,1.5 913.9994374374375u,1.5 914.0004374374374u,0 914.9769774774775u,0 914.9779774774775u,1.5 918.8871376376377u,1.5 918.8881376376377u,0 919.8646776776777u,0 919.8656776776777u,1.5 929.6400780780781u,1.5 929.6410780780781u,0 930.6176181181181u,0 930.6186181181181u,1.5 934.5277782782782u,1.5 934.5287782782782u,0 935.5053183183182u,0 935.5063183183182u,1.5 936.4828583583584u,1.5 936.4838583583584u,0 939.4154784784785u,0 939.4164784784784u,1.5 940.3930185185185u,1.5 940.3940185185185u,0 961.8988993993994u,0 961.8998993993994u,1.5 962.8764394394394u,1.5 962.8774394394394u,0 964.8315195195195u,0 964.8325195195195u,1.5 965.8090595595596u,1.5 965.8100595595596u,0 968.7416796796797u,0 968.7426796796797u,1.5 970.6967597597597u,1.5 970.6977597597597u,0 972.6518398398398u,0 972.6528398398398u,1.5 973.6293798798798u,1.5 973.6303798798798u,0 974.60691991992u,0 974.6079199199199u,1.5 975.58445995996u,1.5 975.58545995996u,0 976.562u,0 976.563u,1.5 977.5395400400402u,1.5 977.5405400400401u,0 978.5170800800801u,0 978.51808008008u,1.5 982.4272402402403u,1.5 982.4282402402403u,0 983.4047802802802u,0 983.4057802802802u,1.5 984.3823203203203u,1.5 984.3833203203203u,0 985.3598603603602u,0 985.3608603603602u,1.5 988.2924804804804u,1.5 988.2934804804804u,0 989.2700205205206u,0 989.2710205205206u,1.5 999.045420920921u,1.5 999.0464209209209u,0 1000.0229609609609u,0 1000.0239609609608u,1.5 1001.000501001001u,1.5 1001.001501001001u,0 1001.9780410410411u,0 1001.9790410410411u,1.5 1011.7534414414415u,1.5 1011.7544414414415u,0 1012.7309814814814u,0 1012.7319814814814u,1.5 1013.7085215215216u,1.5 1013.7095215215215u,0 1014.6860615615615u,0 1014.6870615615614u,1.5 1021.5288418418419u,1.5 1021.5298418418419u,0 1022.5063818818818u,0 1022.5073818818818u,1.5 1023.4839219219219u,1.5 1023.4849219219219u,0 1025.4390020020019u,0 1025.440002002002u,1.5 1026.416542042042u,1.5 1026.4175420420422u,0 1027.394082082082u,0 1027.3950820820821u,1.5 1028.371622122122u,1.5 1028.3726221221223u,0 1029.349162162162u,0 1029.3501621621622u,1.5 1030.3267022022021u,1.5 1030.3277022022023u,0 1031.3042422422423u,0 1031.3052422422425u,1.5 1032.2817822822822u,1.5 1032.2827822822824u,0 1034.2368623623622u,0 1034.2378623623624u,1.5 1035.2144024024024u,1.5 1035.2154024024026u,0 1038.1470225225225u,0 1038.1480225225228u,1.5 1039.1245625625625u,1.5 1039.1255625625627u,0 1063.5630635635634u,0 1063.5640635635636u,1.5 1066.4956836836834u,1.5 1066.4966836836836u,0 1067.4732237237235u,0 1067.4742237237238u,1.5 1085.0689444444445u,1.5 1085.0699444444447u,0 1086.0464844844844u,0 1086.0474844844846u,1.5 1087.0240245245245u,1.5 1087.0250245245247u,0 1088.9791046046046u,0 1088.9801046046048u,1.5 1089.9566446446445u,1.5 1089.9576446446447u,0 1091.9117247247245u,0 1091.9127247247247u,1.5 1092.8892647647647u,1.5 1092.8902647647649u,0 1094.8443448448447u,0 1094.845344844845u,1.5 1095.8218848848846u,1.5 1095.8228848848848u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1120.2603858858856u,1.5 1120.2613858858858u,0 1121.2379259259258u,0 1121.238925925926u,1.5 1122.215465965966u,1.5 1122.216465965966u,0 1123.1930060060058u,0 1123.194006006006u,1.5 1124.170546046046u,1.5 1124.1715460460462u,0 1126.125626126126u,0 1126.1266261261262u,1.5 1127.1031661661661u,1.5 1127.1041661661664u,0 1135.9010265265265u,0 1135.9020265265267u,1.5 1136.8785665665666u,1.5 1136.8795665665668u,0 1137.8561066066065u,0 1137.8571066066067u,1.5 1148.609047047047u,1.5 1148.6100470470471u,0 1149.5865870870869u,0 1149.587587087087u,1.5 1150.564127127127u,1.5 1150.5651271271272u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1174.0250880880878u,1.5 1174.026088088088u,0 1175.9801681681681u,0 1175.9811681681683u,1.5 1176.957708208208u,1.5 1176.9587082082082u,0 1182.8229484484484u,0 1182.8239484484486u,1.5 1183.8004884884883u,1.5 1183.8014884884885u,0 1184.7780285285285u,0 1184.7790285285287u,1.5 1185.7555685685686u,1.5 1185.7565685685688u,0 1186.7331086086085u,0 1186.7341086086087u,1.5 1195.5309689689689u,1.5 1195.531968968969u,0 1196.5085090090088u,0 1196.509509009009u,1.5 1197.486049049049u,1.5 1197.4870490490491u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1214.1042297297297u,1.5 1214.10522972973u,0 1215.0817697697696u,0 1215.0827697697698u,1.5 1217.0368498498497u,1.5 1217.0378498498499u,0 1218.0143898898898u,0 1218.01538988989u,1.5 1218.9919299299297u,1.5 1218.99292992993u,0 1227.7897902902903u,0 1227.7907902902905u,1.5 1229.7448703703703u,1.5 1229.7458703703705u,0 1230.7224104104102u,0 1230.7234104104105u,1.5 1239.5202707707706u,1.5 1239.5212707707708u,0 1241.4753508508506u,0 1241.4763508508508u,1.5 1242.4528908908908u,1.5 1242.453890890891u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1259.0710715715716u,1.5 1259.0720715715718u,0 1261.0261516516516u,0 1261.0271516516518u,1.5 1262.0036916916918u,1.5 1262.004691691692u,0 1264.9363118118117u,0 1264.937311811812u,1.5 1265.9138518518516u,1.5 1265.9148518518518u,0 1268.8464719719718u,0 1268.847471971972u,1.5 1269.8240120120117u,1.5 1269.825012012012u,0 1272.756632132132u,0 1272.7576321321321u,1.5 1282.5320325325324u,1.5 1282.5330325325326u,0 1289.3748128128127u,0 1289.375812812813u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1295.2400530530529u,0 1295.241053053053u,1.5 1299.150213213213u,1.5 1299.1512132132132u,0 1300.127753253253u,0 1300.1287532532533u,1.5 1301.1052932932932u,1.5 1301.1062932932934u,0 1302.0828333333332u,0 1302.0838333333334u,1.5 1303.0603733733733u,1.5 1303.0613733733735u,0 1305.0154534534533u,0 1305.0164534534536u,1.5 1305.9929934934935u,1.5 1305.9939934934937u,0 1314.7908538538536u,0 1314.7918538538538u,1.5 1324.566254254254u,1.5 1324.5672542542543u,0 1325.5437942942942u,0 1325.5447942942944u,1.5 1326.5213343343341u,1.5 1326.5223343343343u,0 1336.2967347347346u,0 1336.2977347347348u,1.5 1337.2742747747748u,1.5 1337.275274774775u,0 1338.251814814815u,0 1338.252814814815u,1.5 1340.2068948948947u,1.5 1340.207894894895u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1350.9598353353351u,1.5 1350.9608353353353u,0 1352.9149154154154u,0 1352.9159154154156u,1.5 1353.8924554554553u,1.5 1353.8934554554555u,0 1361.7127757757758u,0 1361.713775775776u,1.5 1362.690315815816u,1.5 1362.691315815816u,0 1363.6678558558558u,0 1363.668855855856u,1.5 1364.6453958958957u,1.5 1364.646395895896u,0 1365.6229359359356u,0 1365.6239359359358u,1.5 1378.3309564564563u,1.5 1378.3319564564565u,0 1380.2860365365364u,0 1380.2870365365366u,1.5 1381.2635765765765u,1.5 1381.2645765765767u,0 1391.0389769769768u,0 1391.039976976977u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1392.9940570570568u,0 1392.995057057057u,1.5 1393.971597097097u,1.5 1393.9725970970972u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1395.926677177177u,1.5 1395.9276771771772u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1408.6346976976977u,1.5 1408.6356976976979u,0 1409.6122377377376u,0 1409.6132377377378u,1.5 1412.5448578578578u,1.5 1412.545857857858u,0 1413.522397897898u,0 1413.5233978978981u,1.5 1415.4774779779777u,1.5 1415.478477977978u,0 1416.4550180180179u,0 1416.456018018018u,1.5 1417.4325580580578u,1.5 1417.433558058058u,0 1418.410098098098u,0 1418.4110980980981u,1.5 1419.3876381381378u,1.5 1419.388638138138u,0 1436.9833588588588u,0 1436.984358858859u,1.5 1439.915978978979u,1.5 1439.9169789789792u,0 1440.8935190190189u,0 1440.894519019019u,1.5 1441.8710590590588u,1.5 1441.872059059059u,0 1442.848599099099u,0 1442.8495990990991u,1.5 1448.7138393393393u,1.5 1448.7148393393395u,0 1449.6913793793792u,0 1449.6923793793794u,1.5 1463.37693993994u,1.5 1463.3779399399402u,0 1464.35447997998u,0 1464.3554799799801u,1.5 1466.3095600600598u,1.5 1466.31056006006u,0 1467.2871001001u,0 1467.2881001001u,1.5 1468.26464014014u,1.5 1468.2656401401402u,0 1469.24218018018u,0 1469.2431801801802u,1.5 1473.1523403403403u,1.5 1473.1533403403405u,0 1474.1298803803802u,0 1474.1308803803804u,1.5 1476.0849604604603u,1.5 1476.0859604604605u,0 1478.0400405405405u,0 1478.0410405405407u,1.5 1479.0175805805804u,1.5 1479.0185805805806u,0 1482.9277407407408u,0 1482.928740740741u,1.5 1483.9052807807807u,1.5 1483.906280780781u,0 1486.8379009009009u,0 1486.838900900901u,1.5 1487.815440940941u,1.5 1487.8164409409412u,0 1494.658221221221u,0 1494.6592212212213u,1.5 1495.635761261261u,1.5 1495.6367612612612u,0 1497.5908413413413u,0 1497.5918413413415u,1.5 1498.5683813813812u,1.5 1498.5693813813814u,0 1499.5459214214213u,0 1499.5469214214215u,1.5 1500.5234614614612u,1.5 1500.5244614614614u,0 1506.3887017017016u,0 1506.3897017017018u,1.5 1507.3662417417418u,1.5 1507.367241741742u,0 1512.253941941942u,0 1512.2549419419422u,1.5 1513.231481981982u,1.5 1513.2324819819821u,0 1514.209022022022u,0 1514.2100220220223u,1.5 1515.186562062062u,1.5 1515.1875620620622u,0 1521.0518023023021u,0 1521.0528023023023u,1.5 1522.0293423423423u,1.5 1522.0303423423425u,0 1525.9395025025024u,0 1525.9405025025026u,1.5 1528.8721226226226u,1.5 1528.8731226226228u,0 1529.8496626626625u,0 1529.8506626626627u,1.5 1530.8272027027026u,1.5 1530.8282027027028u,0 1531.8047427427427u,0 1531.805742742743u,1.5 1534.7373628628627u,1.5 1534.738362862863u,0 1535.7149029029028u,0 1535.715902902903u,1.5 1537.669982982983u,1.5 1537.670982982983u,0 1538.647523023023u,0 1538.6485230230232u,1.5 1540.6026031031029u,1.5 1540.603603103103u,0 1541.580143143143u,0 1541.5811431431432u,1.5 1561.130943943944u,1.5 1561.1319439439442u,0 1562.108483983984u,0 1562.109483983984u,1.5 1564.063564064064u,1.5 1564.0645640640641u,0 1566.018644144144u,0 1566.0196441441442u,1.5 1566.996184184184u,1.5 1566.997184184184u,0 1583.614364864865u,0 1583.6153648648651u,1.5 1584.5919049049048u,1.5 1584.592904904905u,0 1587.524525025025u,0 1587.5255250250252u,1.5 1589.479605105105u,1.5 1589.4806051051053u,0 1590.457145145145u,0 1590.4581451451452u,1.5 1601.2100855855854u,1.5 1601.2110855855856u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1608.052865865866u,1.5 1608.053865865866u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1619.7833463463462u,0 1619.7843463463464u,1.5 1620.7608863863861u,1.5 1620.7618863863863u,0 1621.7384264264263u,0 1621.7394264264265u,1.5 1622.7159664664664u,1.5 1622.7169664664666u,0 1623.6935065065063u,0 1623.6945065065065u,1.5 1624.6710465465464u,1.5 1624.6720465465467u,0 1625.6485865865864u,0 1625.6495865865866u,1.5 1633.4689069069068u,1.5 1633.469906906907u,0 1634.446446946947u,0 1634.4474469469471u,1.5 1636.401527027027u,1.5 1636.4025270270272u,0 1637.3790670670671u,0 1637.3800670670673u,1.5 1638.356607107107u,1.5 1638.3576071071072u,0 1639.3341471471472u,0 1639.3351471471474u,1.5 1640.311687187187u,1.5 1640.3126871871873u,0 1649.1095475475474u,0 1649.1105475475476u,1.5 1651.0646276276275u,1.5 1651.0656276276277u,0 1652.0421676676676u,0 1652.0431676676678u,1.5 1658.884947947948u,1.5 1658.8859479479481u,0 1659.8624879879878u,0 1659.863487987988u,1.5 1663.7726481481482u,1.5 1663.7736481481484u,0 1674.5255885885883u,0 1674.5265885885885u,1.5 1685.278529029029u,1.5 1685.2795290290292u,0 1686.256069069069u,0 1686.2570690690693u,1.5 1687.233609109109u,1.5 1687.2346091091092u,0 1696.0314694694694u,0 1696.0324694694696u,1.5 1697.9865495495494u,1.5 1697.9875495495496u,0 1698.9640895895895u,0 1698.9650895895898u,1.5 1706.7844099099098u,1.5 1706.78540990991u,0 1707.76194994995u,0 1707.76294994995u,1.5 1708.73948998999u,1.5 1708.7404899899902u,0 1711.67211011011u,0 1711.6731101101102u,1.5 1712.6496501501501u,1.5 1712.6506501501503u,0 1717.5373503503502u,0 1717.5383503503504u,1.5 1718.5148903903903u,1.5 1718.5158903903905u,0 1719.4924304304302u,0 1719.4934304304304u,1.5 1725.3576706706706u,1.5 1725.3586706706708u,0 1726.3352107107105u,0 1726.3362107107107u,1.5 1730.2453708708708u,1.5 1730.246370870871u,0 1731.2229109109107u,0 1731.223910910911u,1.5 1732.2004509509509u,1.5 1732.201450950951u,0 1739.0432312312312u,0 1739.0442312312314u,1.5 1740.0207712712713u,1.5 1740.0217712712715u,0 1740.998311311311u,0 1740.9993113113112u,1.5 1741.9758513513511u,1.5 1741.9768513513513u,0 1742.9533913913913u,0 1742.9543913913915u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1760.549112112112u,0 1760.5501121121122u,1.5 1770.3245125125122u,1.5 1770.3255125125124u,0 1772.2795925925925u,0 1772.2805925925927u,1.5 1773.2571326326324u,1.5 1773.2581326326326u,0 1774.2346726726726u,0 1774.2356726726728u,1.5 1775.2122127127125u,1.5 1775.2132127127127u,0 1782.054992992993u,0 1782.0559929929932u,1.5 1791.8303933933933u,1.5 1791.8313933933935u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1800.6282537537536u,0 1800.6292537537538u,1.5 1801.6057937937937u,1.5 1801.606793793794u,0 1804.5384139139137u,0 1804.539413913914u,1.5 1811.3811941941942u,1.5 1811.3821941941944u,0 1812.3587342342341u,0 1812.3597342342343u,1.5 1813.3362742742743u,1.5 1813.3372742742745u,0 1814.3138143143142u,0 1814.3148143143144u,1.5 1815.2913543543543u,1.5 1815.2923543543545u,0 1823.1116746746745u,0 1823.1126746746747u,1.5 1824.0892147147147u,1.5 1824.0902147147149u,0 1826.0442947947947u,0 1826.045294794795u,1.5 1827.9993748748748u,1.5 1828.000374874875u,0 1828.976914914915u,0 1828.9779149149151u,1.5 1834.842155155155u,1.5 1834.8431551551553u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1851.4603358358356u,0 1851.4613358358358u,1.5 1861.235736236236u,1.5 1861.2367362362363u,0 1862.2132762762762u,0 1862.2142762762765u,1.5 1865.1458963963964u,1.5 1865.1468963963966u,0 1876.8763768768767u,0 1876.877376876877u,1.5 1877.853916916917u,1.5 1877.854916916917u,0 1878.8314569569568u,0 1878.832456956957u,1.5 1880.7865370370369u,1.5 1880.787537037037u,0 1881.764077077077u,0 1881.7650770770772u,1.5 1887.6293173173174u,1.5 1887.6303173173176u,0 1888.6068573573573u,0 1888.6078573573575u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1891.5394774774772u,0 1891.5404774774775u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1895.4496376376374u,1.5 1895.4506376376376u,0 1913.0453583583583u,0 1913.0463583583585u,1.5 1914.0228983983984u,1.5 1914.0238983983986u,0 1915.0004384384383u,0 1915.0014384384385u,1.5 1931.618619119119u,1.5 1931.6196191191193u,0 1932.596159159159u,0 1932.5971591591592u,1.5 1934.551239239239u,1.5 1934.5522392392393u,0 1936.5063193193193u,0 1936.5073193193195u,1.5 1937.4838593593593u,1.5 1937.4848593593595u,0 1938.4613993993994u,0 1938.4623993993996u,1.5 1939.4389394394395u,1.5 1939.4399394394397u,0 1960.94482032032u,0 1960.9458203203203u,1.5 1961.9223603603602u,1.5 1961.9233603603604u,0 1967.7876006006004u,0 1967.7886006006006u,1.5 1969.7426806806807u,1.5 1969.7436806806809u,0 1970.7202207207204u,0 1970.7212207207206u,1.5 1971.6977607607605u,1.5 1971.6987607607607u,0 1972.6753008008006u,0 1972.6763008008008u,1.5 1973.6528408408408u,1.5 1973.653840840841u,0 1974.630380880881u,0 1974.6313808808811u,1.5 1975.6079209209206u,1.5 1975.6089209209208u,0 1976.5854609609607u,0 1976.586460960961u,1.5 1978.540541041041u,1.5 1978.5415410410412u,0 1979.5180810810812u,0 1979.5190810810814u,1.5 1988.3159414414415u,1.5 1988.3169414414417u,0 1989.2934814814816u,0 1989.2944814814819u,1.5 1997.1138018018016u,1.5 1997.1148018018018u,0 1998.0913418418418u,0 1998.092341841842u,1.5 2002.979042042042u,1.5 2002.9800420420422u,0 2003.9565820820822u,0 2003.9575820820824u,1.5 2005.911662162162u,1.5 2005.9126621621622u,0 2006.8892022022021u,0 2006.8902022022023u,1.5 2017.6421426426425u,1.5 2017.6431426426427u,0 2018.6196826826827u,0 2018.6206826826829u,1.5 2020.5747627627625u,1.5 2020.5757627627627u,0 2021.5523028028026u,0 2021.5533028028028u,1.5 2024.4849229229226u,1.5 2024.4859229229228u,0 2025.4624629629627u,0 2025.463462962963u,1.5 2027.417543043043u,1.5 2027.4185430430432u,0 2030.350163163163u,0 2030.3511631631632u,1.5 2031.327703203203u,1.5 2031.3287032032033u,0 2032.3052432432432u,0 2032.3062432432434u,1.5 2033.2827832832834u,1.5 2033.2837832832836u,0 2038.1704834834836u,0 2038.1714834834838u,1.5 2039.1480235235233u,1.5 2039.1490235235235u,0 2058.698824324324u,0 2058.6998243243243u,1.5 2059.676364364364u,1.5 2059.677364364364u,0 2061.6314444444442u,0 2061.6324444444444u,1.5 2062.6089844844846u,1.5 2062.609984484485u,0 2064.5640645645644u,0 2064.5650645645646u,1.5 2065.5416046046043u,1.5 2065.5426046046045u,0 2066.5191446446447u,0 2066.520144644645u,1.5 2068.4742247247245u,1.5 2068.4752247247247u,0 2069.4517647647644u,0 2069.4527647647647u,1.5 2072.384384884885u,1.5 2072.3853848848853u,0 2073.3619249249246u,0 2073.3629249249248u,1.5 2088.025025525525u,1.5 2088.0260255255253u,0 2104.643206206206u,0 2104.644206206206u,1.5 2107.575826326326u,1.5 2107.576826326326u,0 2108.553366366366u,0 2108.554366366366u,1.5 2112.463526526526u,1.5 2112.4645265265262u,0 2113.4410665665664u,0 2113.4420665665666u,1.5 2122.2389269269265u,1.5 2122.2399269269267u,0 2123.216466966967u,0 2123.217466966967u,1.5 2124.194007007007u,1.5 2124.195007007007u,0 2125.171547047047u,0 2125.1725470470474u,1.5 2126.149087087087u,1.5 2126.1500870870873u,0 2136.9020275275275u,0 2136.9030275275277u,1.5 2147.654967967968u,1.5 2147.655967967968u,0 2148.632508008008u,0 2148.633508008008u,1.5 2149.610048048048u,1.5 2149.6110480480484u,0 2161.3405285285285u,0 2161.3415285285287u,1.5 2166.228228728729u,1.5 2166.229228728729u,0 2167.2057687687684u,0 2167.2067687687686u,1.5 2172.093468968969u,1.5 2172.094468968969u,0 2173.071009009009u,0 2173.072009009009u,1.5 2175.026089089089u,1.5 2175.0270890890893u,0 2177.9587092092092u,0 2177.9597092092094u,1.5 2178.936249249249u,1.5 2178.9372492492494u,0 2186.7565695695694u,0 2186.7575695695696u,1.5 2196.53196996997u,1.5 2196.53296996997u,0 2198.48705005005u,0 2198.4880500500503u,1.5 2199.46459009009u,1.5 2199.4655900900902u,0 2201.41967017017u,0 2201.42067017017u,1.5 2202.3972102102102u,1.5 2202.3982102102104u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2219.015390890891u,1.5 2219.016390890891u,0 2229.7683313313314u,0 2229.7693313313316u,1.5 2232.700951451451u,1.5 2232.7019514514514u,0 2233.6784914914915u,0 2233.6794914914917u,1.5 2240.5212717717714u,1.5 2240.5222717717716u,0 2241.4988118118117u,0 2241.499811811812u,1.5 2242.4763518518516u,1.5 2242.477351851852u,0 2250.296672172172u,0 2250.297672172172u,1.5 2258.1169924924925u,1.5 2258.1179924924927u,0 2259.0945325325324u,0 2259.0955325325326u,1.5 2261.0496126126122u,1.5 2261.0506126126124u,0 2262.0271526526526u,0 2262.028152652653u,1.5 2263.0046926926925u,1.5 2263.0056926926927u,0 2270.8250130130127u,0 2270.826013013013u,1.5 2271.802553053053u,1.5 2271.8035530530533u,0 2272.780093093093u,0 2272.781093093093u,1.5 2281.577953453453u,1.5 2281.5789534534533u,0 2291.3533538538536u,0 2291.354353853854u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2294.285973973974u,0 2294.286973973974u,1.5 2304.0613743743743u,1.5 2304.0623743743745u,0 2313.8367747747743u,0 2313.8377747747745u,1.5 2317.746934934935u,1.5 2317.747934934935u,0 2318.724474974975u,0 2318.725474974975u,1.5 2326.5447952952954u,1.5 2326.5457952952956u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2348.050676176176u,1.5 2348.051676176176u,0 2349.028216216216u,0 2349.0292162162164u,1.5 2350.9832962962964u,1.5 2350.9842962962966u,0 2353.915916416416u,0 2353.9169164164164u,1.5 2354.893456456456u,1.5 2354.8944564564563u,0 2360.7586966966965u,0 2360.7596966966967u,1.5 2361.736236736737u,1.5 2361.737236736737u,0 2363.6913168168167u,0 2363.692316816817u,1.5 2364.6688568568566u,1.5 2364.6698568568568u,0 2365.646396896897u,0 2365.647396896897u,1.5 2378.354417417417u,1.5 2378.3554174174174u,0 2379.331957457457u,0 2379.3329574574573u,1.5 2380.3094974974974u,1.5 2380.3104974974976u,0 2388.1298178178176u,0 2388.130817817818u,1.5 2389.1073578578576u,1.5 2389.1083578578578u,0 2393.0175180180177u,0 2393.018518018018u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2394.972598098098u,0 2394.973598098098u,1.5 2395.9501381381383u,1.5 2395.9511381381385u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2398.882758258258u,1.5 2398.8837582582582u,0 2399.8602982982984u,0 2399.8612982982986u,1.5 2408.6581586586585u,1.5 2408.6591586586587u,0 2409.6356986986984u,0 2409.6366986986986u,1.5 2413.5458588588585u,1.5 2413.5468588588587u,0 2430.1640395395393u,0 2430.1650395395395u,1.5 2431.1415795795797u,1.5 2431.14257957958u,0 2433.0966596596595u,0 2433.0976596596597u,1.5 2434.0741996996994u,1.5 2434.0751996996996u,0 2436.0292797797797u,0 2436.03027977978u,1.5 2437.0068198198196u,1.5 2437.00781981982u,0 2438.9618998999u,0 2438.9628998999u,1.5 2463.400400900901u,1.5 2463.401400900901u,0 2465.355480980981u,0 2465.3564809809814u,1.5 2466.3330210210206u,1.5 2466.334021021021u,0 2467.310561061061u,0 2467.311561061061u,1.5 2469.2656411411413u,1.5 2469.2666411411415u,0 2470.243181181181u,0 2470.2441811811814u,1.5 2472.198261261261u,1.5 2472.199261261261u,0 2473.1758013013014u,0 2473.1768013013016u,1.5 2475.1308813813816u,1.5 2475.131881381382u,0 2476.108421421421u,0 2476.1094214214213u,1.5 2477.0859614614615u,1.5 2477.0869614614617u,0 2480.0185815815817u,0 2480.019581581582u,1.5 2480.996121621621u,1.5 2480.9971216216213u,0 2484.9062817817817u,0 2484.907281781782u,1.5 2485.8838218218216u,1.5 2485.884821821822u,0 2487.838901901902u,0 2487.839901901902u,1.5 2488.816441941942u,1.5 2488.817441941942u,0 2494.681682182182u,0 2494.6826821821824u,1.5 2495.659222222222u,1.5 2495.6602222222223u,0 2502.5020025025024u,0 2502.5030025025026u,1.5 2503.4795425425427u,1.5 2503.480542542543u,0 2504.4570825825826u,0 2504.458082582583u,1.5 2505.434622622622u,1.5 2505.4356226226223u,0 2507.3897027027024u,0 2507.3907027027026u,1.5 2508.3672427427427u,1.5 2508.368242742743u,0 2511.2998628628625u,0 2511.3008628628627u,1.5 2512.277402902903u,1.5 2512.278402902903u,0 2513.2549429429428u,0 2513.255942942943u,1.5 2514.232482982983u,1.5 2514.2334829829833u,0 2515.2100230230226u,0 2515.211023023023u,1.5 2516.187563063063u,1.5 2516.188563063063u,0 2522.0528033033033u,0 2522.0538033033035u,1.5 2523.0303433433432u,1.5 2523.0313433433435u,0 2524.0078833833836u,0 2524.008883383384u,1.5 2524.985423423423u,1.5 2524.9864234234233u,0 2526.9405035035034u,0 2526.9415035035036u,1.5 2527.9180435435437u,1.5 2527.919043543544u,0 2528.8955835835836u,0 2528.896583583584u,1.5 2530.8506636636635u,1.5 2530.8516636636637u,0 2531.8282037037034u,0 2531.8292037037036u,1.5 2532.8057437437437u,1.5 2532.806743743744u,0 2533.7832837837836u,0 2533.784283783784u,1.5 2535.7383638638635u,1.5 2535.7393638638637u,0 2536.715903903904u,0 2536.716903903904u,1.5 2540.626064064064u,1.5 2540.627064064064u,0 2541.603604104104u,0 2541.604604104104u,1.5 2563.109484984985u,1.5 2563.1104849849853u,0 2564.0870250250246u,0 2564.0880250250248u,1.5 2566.042105105105u,1.5 2566.043105105105u,0 2568.974725225225u,0 2568.9757252252252u,1.5 2569.952265265265u,1.5 2569.953265265265u,0 2570.9298053053053u,0 2570.9308053053055u,1.5 2571.907345345345u,1.5 2571.9083453453454u,0 2579.7276656656654u,0 2579.7286656656656u,1.5 2580.7052057057053u,1.5 2580.7062057057055u,0 2581.6827457457457u,0 2581.683745745746u,1.5 2582.6602857857856u,1.5 2582.661285785786u,0 2588.5255260260255u,0 2588.5265260260257u,1.5 2590.480606106106u,1.5 2590.481606106106u,0 2591.458146146146u,0 2591.4591461461464u,1.5 2592.435686186186u,1.5 2592.4366861861863u,0 2593.413226226226u,0 2593.414226226226u,1.5 2601.2335465465467u,1.5 2601.234546546547u,0 2602.2110865865866u,0 2602.212086586587u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2607.0987867867866u,1.5 2607.099786786787u,0 2620.784347347347u,0 2620.7853473473474u,1.5 2623.7169674674674u,1.5 2623.7179674674676u,0 2624.6945075075073u,0 2624.6955075075075u,1.5 2625.6720475475477u,1.5 2625.673047547548u,0 2626.6495875875876u,0 2626.650587587588u,1.5 2636.424987987988u,1.5 2636.4259879879883u,0 2638.380068068068u,0 2638.381068068068u,1.5 2639.357608108108u,1.5 2639.358608108108u,0 2648.1554684684684u,0 2648.1564684684686u,1.5 2649.1330085085083u,1.5 2649.1340085085085u,0 2650.1105485485486u,0 2650.111548548549u,1.5 2652.065628628629u,1.5 2652.066628628629u,0 2653.0431686686684u,0 2653.0441686686686u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2673.5715095095093u,0 2673.5725095095095u,1.5 2674.5490495495496u,1.5 2674.55004954955u,0 2676.50412962963u,0 2676.50512962963u,1.5 2686.27953003003u,1.5 2686.28053003003u,0 2687.25707007007u,0 2687.25807007007u,1.5 2688.2346101101098u,1.5 2688.23561011011u,0 2698.0100105105103u,0 2698.0110105105105u,1.5 2698.9875505505506u,1.5 2698.988550550551u,0 2699.9650905905905u,0 2699.9660905905907u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2708.7629509509507u,0 2708.763950950951u,1.5 2709.740490990991u,1.5 2709.741490990991u,0 2716.583271271271u,0 2716.584271271271u,1.5 2718.538351351351u,1.5 2718.5393513513513u,0 2719.5158913913915u,0 2719.5168913913917u,1.5 2721.4709714714713u,1.5 2721.4719714714715u,0 2722.4485115115112u,0 2722.4495115115114u,1.5 2726.3586716716713u,1.5 2726.3596716716715u,0 2727.3362117117117u,0 2727.337211711712u,1.5 2728.3137517517516u,1.5 2728.314751751752u,0 2729.2912917917915u,0 2729.2922917917917u,1.5 2731.2463718718714u,1.5 2731.2473718718716u,0 2735.156532032032u,0 2735.157532032032u,1.5 2736.134072072072u,1.5 2736.135072072072u,0 2739.066692192192u,0 2739.067692192192u,1.5 2740.0442322322324u,1.5 2740.0452322322326u,0 2741.021772272272u,0 2741.022772272272u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2758.617492992993u,0 2758.618492992993u,1.5 2759.595033033033u,1.5 2759.596033033033u,0 2760.572573073073u,0 2760.573573073073u,1.5 2763.505193193193u,1.5 2763.506193193193u,0 2764.4827332332334u,0 2764.4837332332336u,1.5 2768.3928933933935u,1.5 2768.3938933933937u,0 2769.3704334334334u,0 2769.3714334334336u,1.5 2770.3479734734733u,1.5 2770.3489734734735u,0 2771.325513513513u,0 2771.3265135135134u,1.5 2772.3030535535536u,1.5 2772.304053553554u,0 2782.0784539539536u,0 2782.079453953954u,1.5 2790.876314314314u,1.5 2790.8773143143144u,0 2791.853854354354u,0 2791.8548543543543u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2793.8089344344344u,0 2793.8099344344346u,1.5 2794.7864744744743u,1.5 2794.7874744744745u,0 2804.561874874875u,0 2804.562874874875u,1.5 2814.337275275275u,1.5 2814.338275275275u,0 2821.1800555555556u,0 2821.1810555555558u,1.5 2822.1575955955955u,1.5 2822.1585955955957u,0 2828.022835835836u,0 2828.023835835836u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2846.5960965965965u,0 2846.5970965965967u,1.5 2847.573636636637u,1.5 2847.574636636637u,0 2848.5511766766763u,0 2848.5521766766765u,1.5 2849.5287167167166u,1.5 2849.529716716717u,0 2850.5062567567566u,0 2850.5072567567568u,1.5 2851.483796796797u,1.5 2851.484796796797u,0 2852.461336836837u,0 2852.462336836837u,1.5 2861.259197197197u,1.5 2861.260197197197u,0 2862.2367372372373u,0 2862.2377372372375u,1.5 2864.191817317317u,1.5 2864.1928173173173u,0 2876.899837837838u,0 2876.900837837838u,1.5 2877.877377877878u,1.5 2877.8783778778784u,0 2878.8549179179176u,0 2878.855917917918u,1.5 2880.809997997998u,1.5 2880.810997997998u,0 2881.787538038038u,0 2881.788538038038u,1.5 2882.765078078078u,1.5 2882.7660780780784u,0 2883.7426181181177u,0 2883.743618118118u,1.5 2889.607858358358u,1.5 2889.6088583583582u,0 2890.5853983983984u,0 2890.5863983983986u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2897.4281786786787u,0 2897.429178678679u,1.5 2898.4057187187186u,1.5 2898.406718718719u,0 2907.203579079079u,0 2907.2045790790794u,1.5 2908.1811191191186u,1.5 2908.182119119119u,0 2911.1137392392393u,0 2911.1147392392395u,1.5 2912.091279279279u,1.5 2912.0922792792794u,0 2913.068819319319u,0 2913.0698193193193u,1.5 2918.9340595595595u,1.5 2918.9350595595597u,0 2919.9115995995994u,0 2919.9125995995996u,1.5 2928.70945995996u,1.5 2928.71045995996u,0 2929.687u,0 2929.688u,1.5 2933.59716016016u,1.5 2933.59816016016u,0 2934.5747002002u,0 2934.5757002002u,1.5 2935.5522402402403u,1.5 2935.5532402402405u,0 2936.52978028028u,0 2936.5307802802804u,1.5 2937.50732032032u,1.5 2937.5083203203203u,0 2939.4624004004004u,0 2939.4634004004006u,1.5 2940.4399404404403u,1.5 2940.4409404404405u,0 2942.39502052052u,0 2942.3960205205203u,1.5 2943.3725605605605u,1.5 2943.3735605605607u,0 2956.080581081081u,0 2956.0815810810814u,1.5 2957.0581211211206u,1.5 2957.059121121121u,0 2960.968281281281u,0 2960.9692812812814u,1.5 2961.945821321321u,1.5 2961.9468213213213u,0 2962.923361361361u,0 2962.924361361361u,1.5 2964.8784414414413u,1.5 2964.8794414414415u,0 2965.8559814814816u,0 2965.856981481482u,1.5 2966.833521521521u,1.5 2966.8345215215213u,0 2967.8110615615615u,0 2967.8120615615617u,1.5 2968.7886016016014u,1.5 2968.7896016016016u,0 2969.7661416416418u,0 2969.767141641642u,1.5 2970.7436816816817u,1.5 2970.744681681682u,0 2972.6987617617615u,0 2972.6997617617617u,1.5 2974.6538418418418u,1.5 2974.654841841842u,0 2975.631381881882u,0 2975.6323818818823u,1.5 2980.519082082082u,1.5 2980.5200820820824u,0 2981.4966221221216u,0 2981.497622122122u,1.5 2983.451702202202u,1.5 2983.452702202202u,0 2984.4292422422423u,0 2984.4302422422425u,1.5 2986.384322322322u,1.5 2986.3853223223223u,0 2987.361862362362u,0 2987.362862362362u,1.5 2989.3169424424423u,1.5 2989.3179424424425u,0 2990.2944824824826u,0 2990.295482482483u,1.5 2993.2271026026024u,1.5 2993.2281026026026u,0 2994.2046426426427u,0 2994.205642642643u,1.5 2999.0923428428428u,1.5 2999.093342842843u,0 3000.069882882883u,0 3000.0708828828833u,1.5 3003.980043043043u,1.5 3003.9810430430434u,0 3004.957583083083u,0 3004.9585830830833u,1.5 3010.822823323323u,1.5 3010.8238233233233u,0 3011.800363363363u,0 3011.801363363363u,1.5 3014.7329834834836u,1.5 3014.733983483484u,0 3015.710523523523u,0 3015.7115235235233u,1.5 3017.6656036036034u,1.5 3017.6666036036036u,0 3018.6431436436437u,0 3018.644143643644u,1.5 3022.553303803804u,1.5 3022.554303803804u,0 3023.5308438438437u,0 3023.531843843844u,1.5 3026.463463963964u,1.5 3026.464463963964u,0 3027.441004004004u,0 3027.442004004004u,1.5 3028.418544044044u,1.5 3028.4195440440444u,0 3029.396084084084u,0 3029.3970840840843u,1.5 3030.373624124124u,1.5 3030.3746241241242u,0 3032.328704204204u,0 3032.329704204204u,1.5 3033.306244244244u,1.5 3033.3072442442444u,0 3036.238864364364u,0 3036.239864364364u,1.5 3037.2164044044043u,1.5 3037.2174044044045u,0 3039.1714844844846u,0 3039.172484484485u,1.5 3040.149024524524u,1.5 3040.1500245245243u,0 3060.677365365365u,0 3060.678365365365u,1.5 3061.6549054054053u,1.5 3061.6559054054055u,0 3063.6099854854856u,0 3063.610985485486u,1.5 3064.587525525525u,1.5 3064.5885255255253u,0 3065.5650655655654u,0 3065.5660655655656u,1.5 3069.4752257257255u,1.5 3069.4762257257257u,0 3070.4527657657654u,0 3070.4537657657656u,1.5 3074.3629259259255u,1.5 3074.3639259259257u,0 3075.340465965966u,0 3075.341465965966u,1.5 3085.115866366366u,1.5 3085.116866366366u,0 3086.0934064064063u,0 3086.0944064064065u,1.5 3089.026026526526u,1.5 3089.0270265265262u,0 3098.8014269269265u,0 3098.8024269269267u,1.5 3099.778966966967u,1.5 3099.779966966967u,0 3102.711587087087u,0 3102.7125870870873u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3108.576827327327u,1.5 3108.577827327327u,0 3109.554367367367u,0 3109.555367367367u,1.5 3120.307307807808u,1.5 3120.308307807808u,0 3121.2848478478477u,0 3121.285847847848u,1.5 3122.262387887888u,1.5 3122.2633878878883u,0 3132.037788288288u,0 3132.0387882882883u,1.5 3133.0153283283285u,1.5 3133.0163283283287u,0 3134.9704084084083u,0 3134.9714084084085u,1.5 3136.9254884884886u,1.5 3136.9264884884888u,0 3137.9030285285285u,0 3137.9040285285287u,1.5 3145.7233488488487u,1.5 3145.724348848849u,0 3146.700888888889u,0 3146.7018888888892u,1.5 3147.678428928929u,1.5 3147.679428928929u,0 3148.655968968969u,0 3148.656968968969u,1.5 3149.633509009009u,1.5 3149.634509009009u,0 3151.588589089089u,0 3151.5895890890893u,1.5 3152.5661291291294u,1.5 3152.5671291291296u,0 3161.3639894894895u,0 3161.3649894894897u,1.5 3162.3415295295295u,1.5 3162.3425295295297u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3164.2966096096093u,1.5 3164.2976096096095u,0 3165.2741496496496u,0 3165.27514964965u,1.5 3174.0720100100098u,1.5 3174.07301001001u,0 3175.04955005005u,0 3175.0505500500503u,1.5 3176.02709009009u,1.5 3176.0280900900902u,0 3183.8474104104102u,0 3183.8484104104105u,1.5 3184.82495045045u,1.5 3184.8259504504504u,0 3185.8024904904905u,0 3185.8034904904907u,1.5 3186.7800305305304u,1.5 3186.7810305305306u,0 3187.7575705705704u,0 3187.7585705705706u,1.5 3195.577890890891u,1.5 3195.578890890891u,0 3196.555430930931u,0 3196.556430930931u,1.5 3197.532970970971u,1.5 3197.533970970971u,0 3209.263451451451u,0 3209.2644514514514u,1.5 3216.106231731732u,1.5 3216.107231731732u,0 3217.0837717717714u,0 3217.0847717717716u,1.5 3218.0613118118117u,1.5 3218.062311811812u,0 3219.0388518518516u,0 3219.039851851852u,1.5 3220.016391891892u,1.5 3220.017391891892u,0 3229.7917922922925u,0 3229.7927922922927u,1.5 3238.5896526526526u,1.5 3238.590652652653u,0 3240.544732732733u,0 3240.545732732733u,1.5 3241.5222727727723u,1.5 3241.5232727727725u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3261.0730735735733u,1.5 3261.0740735735735u,0 3262.050613613613u,0 3262.0516136136134u,1.5 3263.0281536536536u,1.5 3263.029153653654u,0 3269.870933933934u,0 3269.871933933934u,1.5 3270.848473973974u,1.5 3270.849473973974u,0 3271.8260140140137u,0 3271.827014014014u,1.5 3272.803554054054u,1.5 3272.8045540540543u,0 3273.781094094094u,0 3273.782094094094u,1.5 3280.6238743743743u,1.5 3280.6248743743745u,0 3281.601414414414u,0 3281.6024144144144u,1.5 3283.5564944944945u,1.5 3283.5574944944947u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3301.152215215215u,1.5 3301.1532152152154u,0 3302.129755255255u,0 3302.1307552552553u,1.5 3303.1072952952954u,1.5 3303.1082952952956u,0 3306.039915415415u,0 3306.0409154154154u,1.5 3307.017455455455u,1.5 3307.0184554554553u,0 3312.8826956956955u,0 3312.8836956956957u,1.5 3314.8377757757753u,1.5 3314.8387757757755u,0 3315.8153158158157u,0 3315.816315815816u,1.5 3317.770395895896u,1.5 3317.771395895896u,0 3318.747935935936u,0 3318.748935935936u,1.5 3325.590716216216u,1.5 3325.5917162162164u,0 3326.568256256256u,0 3326.5692562562563u,1.5 3327.5457962962964u,1.5 3327.5467962962966u,0 3328.5233363363363u,0 3328.5243363363365u,1.5 3329.5008763763763u,1.5 3329.5018763763765u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3337.3211966966965u,1.5 3337.3221966966967u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3350.029217217217u,1.5 3350.0302172172173u,0 3351.006757257257u,0 3351.0077572572573u,1.5 3351.9842972972974u,1.5 3351.9852972972976u,0 3361.7596976976974u,0 3361.7606976976977u,1.5 3363.7147777777773u,1.5 3363.7157777777775u,0 3364.6923178178176u,0 3364.693317817818u,1.5 3379.355418418418u,1.5 3379.3564184184183u,0 3382.2880385385383u,0 3382.2890385385385u,1.5 3383.2655785785787u,1.5 3383.266578578579u,0 3388.1532787787787u,0 3388.154278778779u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.0185190190186u,1.5 3394.019519019019u,0 3394.996059059059u,0 3394.997059059059u,1.5 3398.906219219219u,1.5 3398.9072192192193u,0 3399.883759259259u,0 3399.884759259259u,1.5 3408.681619619619u,1.5 3408.6826196196193u,0 3409.6591596596595u,0 3409.6601596596597u,1.5 3410.6366996996994u,1.5 3410.6376996996996u,0 3411.61423973974u,0 3411.61523973974u,1.5 3412.5917797797797u,1.5 3412.59277977978u,0 3414.5468598598595u,0 3414.5478598598597u,1.5 3415.5243998999u,1.5 3415.5253998999u,0 3433.12012062062u,0 3433.1211206206203u,1.5 3435.0752007007004u,1.5 3435.0762007007006u,0 3437.0302807807807u,0 3437.031280780781u,1.5 3438.0078208208206u,1.5 3438.008820820821u,0 3438.9853608608605u,0 3438.9863608608607u,1.5 3460.4912417417418u,1.5 3460.492241741742u,0 3461.4687817817817u,0 3461.469781781782u,1.5 3465.378941941942u,1.5 3465.379941941942u,0 3466.356481981982u,0 3466.3574819819823u,1.5 3467.3340220220216u,1.5 3467.335022022022u,0 3468.311562062062u,0 3468.312562062062u,1.5 3469.289102102102u,1.5 3469.290102102102u,0 3470.2666421421422u,0 3470.2676421421424u,1.5 3472.221722222222u,1.5 3472.2227222222223u,0 3473.199262262262u,0 3473.200262262262u,1.5 3474.1768023023023u,1.5 3474.1778023023026u,0 3475.1543423423423u,0 3475.1553423423425u,1.5 3476.1318823823826u,1.5 3476.132882382383u,0 3478.0869624624625u,0 3478.0879624624627u,1.5 3479.0645025025024u,1.5 3479.0655025025026u,0 3481.0195825825826u,0 3481.020582582583u,1.5 3481.997122622622u,1.5 3481.9981226226223u,0 3482.9746626626625u,0 3482.9756626626627u,1.5 3483.9522027027024u,1.5 3483.9532027027026u,0 3493.727603103103u,0 3493.728603103103u,1.5 3494.7051431431432u,1.5 3494.7061431431434u,0 3501.547923423423u,0 3501.5489234234233u,1.5 3502.5254634634634u,1.5 3502.5264634634636u,0 3521.098724224224u,0 3521.0997242242242u,1.5 3522.076264264264u,1.5 3522.077264264264u,0 3525.0088843843846u,0 3525.009884384385u,1.5 3526.9639644644644u,1.5 3526.9649644644646u,0 3527.9415045045043u,0 3527.9425045045045u,1.5 3529.8965845845846u,1.5 3529.897584584585u,0 3530.8741246246245u,0 3530.8751246246247u,1.5 3531.8516646646644u,1.5 3531.8526646646646u,0 3533.8067447447447u,0 3533.807744744745u,1.5 3535.7618248248245u,1.5 3535.7628248248247u,0 3536.7393648648645u,0 3536.7403648648647u,1.5 3537.716904904905u,1.5 3537.717904904905u,0 3538.6944449449447u,0 3538.695444944945u,1.5 3540.6495250250246u,1.5 3540.6505250250248u,0 3541.627065065065u,0 3541.628065065065u,1.5 3561.1778658658654u,1.5 3561.1788658658656u,0 3562.155405905906u,0 3562.156405905906u,1.5 3564.110485985986u,1.5 3564.1114859859863u,0 3565.0880260260255u,0 3565.0890260260257u,1.5 3566.065566066066u,1.5 3566.066566066066u,0 3568.998186186186u,0 3568.9991861861863u,1.5 3569.975726226226u,1.5 3569.976726226226u,0 3583.6612867867866u,0 3583.662286786787u,1.5 3584.6388268268265u,1.5 3584.6398268268267u,0 3586.593906906907u,0 3586.594906906907u,1.5 3588.548986986987u,1.5 3588.5499869869873u,0 3589.5265270270265u,0 3589.5275270270267u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3609.0773278278275u,1.5 3609.0783278278277u,0 3618.852728228228u,0 3618.853728228228u,1.5 3619.830268268268u,1.5 3619.831268268268u,0 3621.785348348348u,0 3621.7863483483484u,1.5 3622.7628883883885u,1.5 3622.7638883883888u,0 3623.740428428428u,0 3623.741428428428u,1.5 3636.4484489489487u,1.5 3636.449448948949u,0 3638.403529029029u,0 3638.404529029029u,1.5 3639.381069069069u,1.5 3639.382069069069u,0 3650.1340095095093u,0 3650.1350095095095u,1.5 3651.1115495495496u,1.5 3651.11254954955u,0 3652.0890895895895u,0 3652.0900895895898u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3669.6848103103102u,0 3669.6858103103104u,1.5 3670.66235035035u,1.5 3670.6633503503504u,0 3675.5500505505506u,0 3675.551050550551u,1.5 3676.5275905905905u,1.5 3676.5285905905907u,0 3677.505130630631u,0 3677.506130630631u,1.5 3681.4152907907906u,1.5 3681.4162907907908u,0 3682.392830830831u,0 3682.393830830831u,1.5 3685.3254509509507u,1.5 3685.326450950951u,0 3686.302990990991u,0 3686.303990990991u,1.5 3687.280531031031u,1.5 3687.281531031031u,0 3697.0559314314314u,0 3697.0569314314316u,1.5 3698.0334714714713u,1.5 3698.0344714714715u,0 3699.0110115115112u,0 3699.0120115115114u,1.5 3704.8762517517516u,1.5 3704.877251751752u,0 3705.8537917917915u,0 3705.8547917917917u,1.5 3707.8088718718714u,1.5 3707.8098718718716u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3718.561812312312u,0 3718.5628123123124u,1.5 3719.539352352352u,1.5 3719.5403523523523u,0 3720.5168923923925u,0 3720.5178923923927u,1.5 3728.3372127127127u,1.5 3728.338212712713u,0 3729.3147527527526u,0 3729.315752752753u,1.5 3730.292292792793u,1.5 3730.293292792793u,0 3733.2249129129127u,0 3733.225912912913u,1.5 3734.2024529529526u,1.5 3734.203452952953u,0 3740.067693193193u,0 3740.068693193193u,1.5 3746.9104734734733u,1.5 3746.9114734734735u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3758.6409539539536u,0 3758.641953953954u,1.5 3759.618493993994u,1.5 3759.619493993994u,0 3760.596034034034u,0 3760.597034034034u,1.5 3762.5511141141137u,1.5 3762.552114114114u,0 3763.528654154154u,0 3763.5296541541543u,1.5 3770.3714344344344u,1.5 3770.3724344344346u,0 3780.146834834835u,0 3780.147834834835u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3800.6751756756753u,0 3800.6761756756755u,1.5 3801.6527157157157u,1.5 3801.653715715716u,0 3804.585335835836u,0 3804.586335835836u,1.5 3815.338276276276u,1.5 3815.339276276276u,0 3829.023836836837u,0 3829.024836836837u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3851.5072577577575u,0 3851.5082577577577u,1.5 3862.260198198198u,1.5 3862.261198198198u,0 3864.2152782782778u,0 3864.216278278278u,1.5 3865.192818318318u,1.5 3865.1938183183183u,0 3873.013138638639u,0 3873.014138638639u,1.5 3873.9906786786783u,1.5 3873.9916786786785u,0 3877.900838838839u,0 3877.901838838839u,1.5 3878.878378878879u,1.5 3878.8793788788794u,0 3879.8559189189186u,0 3879.856918918919u,1.5 3889.631319319319u,1.5 3889.6323193193193u,0 3890.608859359359u,0 3890.6098593593592u,1.5 3892.5639394394393u,1.5 3892.5649394394395u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3907.22704004004u,0 3907.22804004004u,1.5 3908.20458008008u,1.5 3908.2055800800804u,0 3909.1821201201196u,0 3909.18312012012u,1.5 3910.1596601601605u,1.5 3910.1606601601607u,0 3913.09228028028u,0 3913.0932802802804u,1.5 3929.710460960961u,1.5 3929.711460960961u,0 3930.688001001001u,0 3930.689001001001u,1.5 3931.665541041041u,1.5 3931.666541041041u,0 3932.643081081081u,0 3932.6440810810814u,1.5 3934.5981611611614u,1.5 3934.5991611611616u,0 3935.575701201201u,0 3935.576701201201u,1.5 3937.530781281281u,1.5 3937.5317812812814u,0 3958.0591221221216u,0 3958.060122122122u,1.5 3959.0366621621624u,1.5 3959.0376621621626u,0 3964.9019024024024u,0 3964.9029024024026u,1.5 3965.879442442442u,1.5 3965.880442442442u,0 3967.834522522522u,0 3967.8355225225223u,1.5 3969.7896026026024u,1.5 3969.7906026026026u,0 3970.7671426426423u,0 3970.7681426426425u,1.5 3971.7446826826827u,1.5 3971.745682682683u,0 3972.7222227227226u,0 3972.7232227227228u,1.5 3974.677302802803u,1.5 3974.678302802803u,0 3976.632382882883u,0 3976.6333828828833u,1.5 3977.6099229229226u,1.5 3977.610922922923u,0 3978.5874629629634u,0 3978.5884629629636u,1.5 3985.430243243243u,1.5 3985.431243243243u,0 3986.407783283283u,0 3986.4087832832834u,1.5 3990.317943443443u,1.5 3990.318943443443u,0 3991.2954834834836u,0 3991.296483483484u,1.5 3994.2281036036034u,1.5 3994.2291036036036u,0 3995.2056436436433u,0 3995.2066436436435u,1.5 3998.138263763764u,1.5 3998.139263763764u,0 3999.115803803804u,0 3999.116803803804u,1.5 4004.9810440440438u,1.5 4004.982044044044u,0 4005.958584084084u,0 4005.9595840840843u,1.5 4010.846284284284u,1.5 4010.8472842842843u,0 4011.823824324324u,0 4011.8248243243243u,1.5 4012.8013643643644u,1.5 4012.8023643643646u,0 4013.7789044044043u,0 4013.7799044044045u,1.5 4018.6666046046043u,1.5 4018.6676046046045u,0 4019.6441446446443u,0 4019.6451446446445u,1.5 4023.554304804805u,1.5 4023.555304804805u,0 4024.5318448448443u,0 4024.5328448448445u,1.5 4025.509384884885u,1.5 4025.5103848848853u,0 4026.4869249249246u,0 4026.4879249249248u,1.5 4027.4644649649654u,1.5 4027.4654649649656u,0 4028.442005005005u,0 4028.443005005005u,1.5 4029.4195450450447u,1.5 4029.420545045045u,0 4031.374625125125u,0 4031.375625125125u,1.5 4032.3521651651654u,1.5 4032.3531651651656u,0 4033.329705205205u,0 4033.330705205205u,1.5 4035.284785285285u,1.5 4035.2857852852853u,0 4064.6109864864866u,0 4064.611986486487u,1.5 4068.5211466466462u,1.5 4068.5221466466464u,0 4069.4986866866866u,0 4069.499686686687u,1.5 4070.4762267267265u,1.5 4070.4772267267267u,0 4071.453766766767u,0 4071.454766766767u,1.5 4078.2965470470467u,1.5 4078.297547047047u,0 4079.274087087087u,0 4079.2750870870873u,1.5 4081.2291671671674u,1.5 4081.2301671671676u,0 4082.206707207207u,0 4082.207707207207u,1.5 4087.0944074074073u,1.5 4087.0954074074075u,0 4089.0494874874876u,0 4089.0504874874878u,1.5 4090.027027527527u,1.5 4090.0280275275272u,0 4093.9371876876876u,0 4093.938187687688u,1.5 4094.9147277277275u,1.5 4094.9157277277277u,0 4103.7125880880885u,0 4103.713588088089u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4106.645208208208u,0 4106.646208208208u,1.5 4120.330768768769u,1.5 4120.3317687687695u,0 4121.308308808809u,0 4121.309308808809u,1.5 4122.285848848848u,1.5 4122.286848848848u,0 4124.240928928929u,0 4124.241928928929u,1.5 4125.218468968969u,1.5 4125.2194689689695u,0 4131.083709209209u,0 4131.084709209209u,1.5 4132.061249249249u,1.5 4132.062249249249u,0 4136.948949449449u,0 4136.949949449449u,1.5 4138.904029529529u,1.5 4138.905029529529u,0 4139.881569569569u,0 4139.88256956957u,1.5 4148.67942992993u,1.5 4148.68042992993u,0 4149.65696996997u,0 4149.6579699699705u,1.5 4150.63451001001u,1.5 4150.63551001001u,0 4160.40991041041u,0 4160.41091041041u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4162.3649904904905u,0 4162.365990490491u,1.5 4164.32007057057u,1.5 4164.321070570571u,0 4165.297610610611u,0 4165.298610610611u,1.5 4172.140390890891u,1.5 4172.141390890891u,0 4173.117930930931u,0 4173.118930930931u,1.5 4174.095470970971u,1.5 4174.0964709709715u,0 4185.825951451451u,0 4185.826951451451u,1.5 4186.8034914914915u,1.5 4186.804491491492u,0 4187.781031531531u,0 4187.782031531531u,1.5 4193.646271771772u,1.5 4193.6472717717725u,0 4194.623811811812u,0 4194.624811811812u,1.5 4197.556431931932u,1.5 4197.557431931932u,0 4198.533971971972u,0 4198.5349719719725u,1.5 4199.511512012012u,1.5 4199.512512012012u,0 4206.3542922922925u,0 4206.355292292293u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4210.264452452452u,1.5 4210.265452452452u,0 4211.2419924924925u,0 4211.242992492493u,1.5 4217.107232732732u,1.5 4217.108232732732u,0 4218.084772772773u,0 4218.085772772773u,1.5 4219.062312812813u,1.5 4219.063312812813u,0 4228.837713213213u,0 4228.838713213213u,1.5 4230.7927932932935u,1.5 4230.793793293294u,0 4231.770333333333u,0 4231.771333333333u,1.5 4237.635573573573u,1.5 4237.6365735735735u,0 4238.613113613614u,0 4238.614113613614u,1.5 4240.5681936936935u,1.5 4240.569193693694u,0 4243.500813813814u,0 4243.501813813814u,1.5 4244.478353853853u,1.5 4244.479353853853u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4261.096534534534u,1.5 4261.097534534534u,0 4263.051614614615u,0 4263.052614614615u,1.5 4264.029154654655u,1.5 4264.030154654655u,0 4266.961774774775u,0 4266.962774774775u,1.5 4267.939314814815u,1.5 4267.940314814815u,0 4271.849474974975u,0 4271.850474974975u,1.5 4279.669795295295u,1.5 4279.670795295296u,0 4280.647335335335u,0 4280.648335335335u,1.5 4281.624875375375u,1.5 4281.6258753753755u,0 4293.355355855856u,0 4293.356355855856u,1.5 4301.175676176176u,1.5 4301.176676176176u,0 4302.153216216216u,0 4302.154216216216u,1.5 4303.130756256257u,1.5 4303.131756256257u,0 4315.838776776777u,0 4315.839776776777u,1.5 4316.816316816817u,1.5 4316.817316816817u,0 4317.793856856857u,0 4317.794856856857u,1.5 4325.614177177177u,1.5 4325.615177177177u,0 4326.591717217217u,0 4326.592717217217u,1.5 4327.569257257258u,1.5 4327.570257257258u,0 4328.546797297297u,0 4328.547797297298u,1.5 4329.524337337337u,1.5 4329.525337337337u,0 4334.412037537537u,0 4334.413037537537u,1.5 4335.389577577577u,1.5 4335.3905775775775u,0 4338.322197697697u,0 4338.323197697698u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4351.030218218218u,1.5 4351.031218218218u,0 4352.007758258259u,0 4352.008758258259u,1.5 4352.985298298298u,1.5 4352.986298298299u,0 4360.805618618619u,0 4360.806618618619u,1.5 4361.783158658659u,1.5 4361.784158658659u,0 4363.738238738738u,0 4363.739238738738u,1.5 4365.693318818819u,1.5 4365.694318818819u,0 4366.670858858859u,0 4366.671858858859u,1.5 4376.44625925926u,1.5 4376.44725925926u,0 4377.423799299299u,0 4377.4247992993u,1.5 4379.378879379379u,1.5 4379.379879379379u,0 4392.086899899899u,0 4392.0878998999u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.01952002002u,1.5 4395.02052002002u,0 4396.9746001001u,0 4396.975600100101u,1.5 4407.72754054054u,1.5 4407.72854054054u,0 4408.70508058058u,0 4408.70608058058u,1.5 4409.682620620621u,1.5 4409.683620620621u,0 4410.660160660661u,0 4410.661160660661u,1.5 4412.61524074074u,1.5 4412.61624074074u,0 4414.570320820821u,0 4414.571320820821u,1.5 4415.547860860861u,1.5 4415.548860860861u,0 4430.210961461462u,0 4430.211961461462u,1.5 4431.188501501501u,1.5 4431.189501501502u,0 4432.166041541541u,0 4432.167041541541u,1.5 4434.121121621622u,1.5 4434.122121621622u,0 4435.098661661662u,0 4435.099661661662u,1.5 4436.076201701701u,1.5 4436.077201701702u,0 4437.053741741741u,0 4437.054741741741u,1.5 4439.008821821822u,1.5 4439.009821821822u,0 4439.986361861862u,0 4439.987361861862u,1.5 4440.963901901901u,1.5 4440.964901901902u,0 4441.941441941942u,0 4441.942441941942u,1.5 4457.582082582582u,1.5 4457.583082582582u,0 4458.559622622623u,0 4458.560622622623u,1.5 4459.537162662663u,1.5 4459.538162662663u,0 4460.514702702702u,0 4460.515702702703u,1.5 4467.357482982983u,1.5 4467.358482982983u,0 4468.335023023023u,0 4468.336023023023u,1.5 4469.312563063063u,1.5 4469.313563063063u,0 4471.267643143143u,0 4471.268643143143u,1.5 4472.245183183183u,1.5 4472.246183183183u,0 4473.222723223223u,0 4473.223723223223u,1.5 4474.200263263264u,1.5 4474.201263263264u,0 4475.177803303303u,0 4475.1788033033035u,1.5 4476.155343343343u,1.5 4476.156343343343u,0 4478.1104234234235u,0 4478.111423423424u,1.5 4479.087963463464u,1.5 4479.088963463464u,0 4482.9981236236235u,0 4482.999123623624u,1.5 4483.975663663664u,1.5 4483.976663663664u,0 4484.953203703703u,0 4484.954203703704u,1.5 4485.930743743743u,1.5 4485.931743743743u,0 4491.795983983984u,0 4491.796983983984u,1.5 4492.773524024024u,1.5 4492.774524024024u,0 4494.728604104104u,0 4494.7296041041045u,1.5 4495.706144144144u,1.5 4495.707144144144u,0 4503.526464464465u,0 4503.527464464465u,1.5 4504.504004504504u,1.5 4504.5050045045045u,0 4506.459084584585u,0 4506.460084584585u,1.5 4507.4366246246245u,1.5 4507.437624624625u,0 4510.369244744744u,0 4510.370244744744u,1.5 4511.346784784785u,1.5 4511.347784784785u,0 4514.279404904904u,0 4514.280404904905u,1.5 4515.256944944945u,1.5 4515.257944944945u,0 4519.167105105105u,0 4519.1681051051055u,1.5 4520.144645145145u,1.5 4520.145645145145u,0 4522.099725225225u,0 4522.100725225225u,1.5 4523.077265265266u,1.5 4523.078265265266u,0 4525.032345345345u,0 4525.033345345345u,1.5 4526.9874254254255u,1.5 4526.988425425426u,0 4528.942505505505u,0 4528.9435055055055u,1.5 4529.920045545545u,1.5 4529.921045545545u,0 4531.8751256256255u,0 4531.876125625626u,1.5 4536.7628258258255u,1.5 4536.763825825826u,0 4537.740365865866u,0 4537.741365865866u,1.5 4539.695445945946u,1.5 4539.696445945946u,0 4540.672985985986u,0 4540.673985985986u,1.5 4542.628066066066u,1.5 4542.629066066066u,0 4543.605606106106u,0 4543.6066061061065u,1.5 4562.178866866867u,1.5 4562.179866866867u,0 4563.156406906906u,0 4563.1574069069065u,1.5 4565.111486986987u,1.5 4565.112486986987u,0 4569.021647147147u,0 4569.022647147147u,1.5 4569.999187187187u,1.5 4570.000187187187u,0 4584.662287787788u,0 4584.663287787788u,1.5 4585.6398278278275u,1.5 4585.640827827828u,0 4586.617367867868u,0 4586.618367867868u,1.5 4587.594907907907u,1.5 4587.5959079079075u,0 4588.572447947948u,0 4588.573447947948u,1.5 4590.5275280280275u,1.5 4590.528528028028u,0 4591.505068068068u,0 4591.506068068068u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4607.145708708708u,0 4607.1467087087085u,1.5 4608.123248748749u,1.5 4608.124248748749u,0 4620.83126926927u,0 4620.83226926927u,1.5 4622.786349349349u,1.5 4622.787349349349u,0 4623.763889389389u,0 4623.764889389389u,1.5 4634.5168298298295u,1.5 4634.51782982983u,0 4635.49436986987u,0 4635.49536986987u,1.5 4637.44944994995u,1.5 4637.45044994995u,0 4640.38207007007u,0 4640.38307007007u,1.5 4641.35961011011u,1.5 4641.36061011011u,0 4649.17993043043u,0 4649.180930430431u,1.5 4651.13501051051u,1.5 4651.1360105105105u,0 4652.11255055055u,0 4652.11355055055u,1.5 4653.090090590591u,1.5 4653.091090590591u,0 4654.06763063063u,0 4654.068630630631u,1.5 4659.932870870871u,1.5 4659.933870870871u,0 4660.91041091091u,0 4660.9114109109105u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4666.775651151151u,0 4666.776651151151u,1.5 4667.753191191191u,1.5 4667.754191191191u,0 4671.663351351351u,0 4671.664351351351u,1.5 4672.640891391391u,1.5 4672.641891391391u,0 4673.618431431431u,0 4673.619431431432u,1.5 4685.348911911911u,1.5 4685.3499119119115u,0 4686.326451951952u,0 4686.327451951952u,1.5 4687.303991991992u,1.5 4687.304991991992u,0 4688.2815320320315u,0 4688.282532032032u,1.5 4689.259072072072u,1.5 4689.260072072072u,0 4697.079392392392u,0 4697.080392392392u,1.5 4698.056932432432u,1.5 4698.057932432433u,0 4699.034472472473u,0 4699.035472472473u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4709.787412912912u,1.5 4709.7884129129125u,0 4718.585273273274u,0 4718.586273273274u,1.5 4720.540353353353u,1.5 4720.541353353353u,0 4721.517893393393u,0 4721.518893393393u,1.5 4726.405593593594u,1.5 4726.406593593594u,0 4727.383133633633u,0 4727.384133633634u,1.5 4729.338213713713u,1.5 4729.339213713713u,0 4740.091154154154u,0 4740.092154154154u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4760.619494994995u,0 4760.620494994995u,1.5 4761.597035035034u,1.5 4761.598035035035u,0 4762.574575075075u,0 4762.575575075075u,1.5 4770.394895395395u,1.5 4770.395895395395u,0 4772.349975475476u,0 4772.350975475476u,1.5 4773.327515515515u,1.5 4773.328515515515u,0 4777.237675675676u,0 4777.238675675676u,1.5 4778.215215715715u,1.5 4778.216215715715u,0 4781.147835835835u,0 4781.148835835836u,1.5 4784.0804559559565u,1.5 4784.081455955957u,0 4785.057995995996u,0 4785.058995995996u,1.5 4792.878316316316u,1.5 4792.879316316316u,0 4795.810936436436u,0 4795.811936436437u,1.5 4796.788476476477u,1.5 4796.789476476477u,0 4804.608796796797u,0 4804.609796796797u,1.5 4815.361737237236u,1.5 4815.362737237237u,0 4816.339277277278u,0 4816.340277277278u,1.5 4817.316817317317u,1.5 4817.317817317317u,0 4823.1820575575575u,0 4823.183057557558u,1.5 4824.159597597598u,1.5 4824.160597597598u,0 4825.137137637637u,0 4825.138137637638u,1.5 4826.114677677678u,1.5 4826.115677677678u,0 4827.092217717717u,0 4827.093217717717u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4849.575638638638u,0 4849.5766386386385u,1.5 4850.553178678679u,1.5 4850.554178678679u,0 4851.530718718718u,0 4851.531718718718u,1.5 4852.508258758759u,1.5 4852.50925875876u,0 4853.485798798799u,0 4853.486798798799u,1.5 4865.21627927928u,1.5 4865.21727927928u,0 4876.94675975976u,0 4876.947759759761u,1.5 4877.9242997998u,1.5 4877.9252997998u,0 4878.901839839839u,0 4878.9028398398395u,1.5 4879.87937987988u,1.5 4879.88037987988u,0 4880.85691991992u,0 4880.85791991992u,1.5 4882.812u,1.5 4882.813u,0 4883.789540040039u,0 4883.79054004004u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4895.52002052052u,0 4895.52102052052u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4907.250501001001u,0 4907.251501001001u,1.5 4908.22804104104u,1.5 4908.229041041041u,0 4911.160661161161u,0 4911.161661161162u,1.5 4912.138201201201u,1.5 4912.139201201201u,0 4914.093281281282u,0 4914.094281281282u,1.5 4917.025901401401u,1.5 4917.026901401401u,0 4918.003441441441u,0 4918.0044414414415u,1.5 4930.711461961962u,1.5 4930.712461961963u,0 4931.689002002002u,0 4931.690002002002u,1.5 4933.644082082082u,1.5 4933.645082082082u,0 4934.621622122122u,0 4934.622622122122u,1.5 4935.599162162162u,1.5 4935.600162162163u,0 4936.576702202202u,0 4936.577702202202u,1.5 4937.554242242241u,1.5 4937.555242242242u,0 4939.509322322322u,0 4939.510322322322u,1.5 4940.486862362362u,1.5 4940.487862362363u,0 4964.925363363363u,0 4964.926363363364u,1.5 4965.902903403403u,1.5 4965.903903403403u,0 4969.813063563563u,0 4969.814063563564u,1.5 4970.790603603604u,1.5 4970.791603603604u,0 4971.768143643643u,0 4971.7691436436435u,1.5 4972.745683683684u,1.5 4972.746683683684u,0 4973.723223723723u,0 4973.724223723723u,1.5 4974.700763763764u,1.5 4974.701763763765u,0 4976.655843843843u,0 4976.6568438438435u,1.5 4977.633383883884u,1.5 4977.634383883884u,0 4978.610923923924u,0 4978.611923923924u,1.5 4983.498624124124u,1.5 4983.499624124124u,0 4984.476164164164u,0 4984.477164164165u,1.5 4988.386324324324u,1.5 4988.387324324324u,0 4989.363864364364u,0 4989.364864364365u,1.5 5003.049424924925u,1.5 5003.050424924925u,0 5004.026964964965u,0 5004.027964964966u,1.5 5005.982045045044u,1.5 5005.9830450450445u,0 5006.959585085086u,0 5006.960585085086u,1.5 5014.779905405405u,1.5 5014.780905405405u,0 5015.757445445445u,0 5015.758445445445u,1.5 5017.712525525525u,1.5 5017.713525525525u,0 5018.690065565565u,0 5018.691065565566u,1.5 5020.645145645645u,1.5 5020.646145645645u,0 5021.622685685686u,0 5021.623685685686u,1.5 5022.600225725725u,1.5 5022.601225725725u,0 5024.555305805806u,0 5024.556305805806u,1.5 5025.532845845845u,1.5 5025.5338458458455u,0 5026.510385885886u,0 5026.511385885886u,1.5 5028.465465965966u,1.5 5028.466465965967u,0 5029.443006006006u,0 5029.444006006006u,1.5 5031.398086086087u,1.5 5031.399086086087u,0 5033.353166166166u,0 5033.354166166167u,1.5 5034.330706206206u,1.5 5034.331706206206u,0 5042.151026526526u,0 5042.152026526526u,1.5 5043.128566566566u,1.5 5043.129566566567u,0 5055.8365870870875u,0 5055.837587087088u,1.5 5056.814127127127u,1.5 5056.815127127127u,0 5059.746747247247u,0 5059.747747247247u,1.5 5060.724287287288u,1.5 5060.725287287288u,0 5061.701827327327u,0 5061.702827327327u,1.5 5062.679367367367u,1.5 5062.680367367368u,0 5063.656907407407u,0 5063.657907407407u,1.5 5065.611987487488u,1.5 5065.612987487488u,0 5066.589527527527u,0 5066.590527527527u,1.5 5067.567067567567u,1.5 5067.568067567568u,0 5068.544607607608u,0 5068.545607607608u,1.5 5071.477227727727u,1.5 5071.478227727727u,0 5072.454767767768u,0 5072.4557677677685u,1.5 5084.185248248248u,1.5 5084.186248248248u,0 5085.1627882882885u,0 5085.163788288289u,1.5 5087.117868368368u,1.5 5087.118868368369u,0 5088.095408408408u,0 5088.096408408408u,1.5 5089.072948448448u,1.5 5089.073948448448u,0 5092.983108608609u,0 5092.984108608609u,1.5 5093.960648648648u,1.5 5093.961648648648u,0 5095.915728728728u,0 5095.916728728728u,1.5 5096.893268768769u,1.5 5096.8942687687695u,0 5103.736049049048u,0 5103.737049049048u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5108.623749249249u,0 5108.624749249249u,1.5 5117.42160960961u,1.5 5117.42260960961u,0 5118.399149649649u,0 5118.400149649649u,1.5 5121.33176976977u,1.5 5121.3327697697705u,0 5122.30930980981u,0 5122.31030980981u,1.5 5123.286849849849u,1.5 5123.287849849849u,0 5134.0397902902905u,0 5134.040790290291u,1.5 5135.01733033033u,1.5 5135.01833033033u,0 5136.97241041041u,0 5136.97341041041u,1.5 5137.94995045045u,1.5 5137.95095045045u,0 5138.9274904904905u,0 5138.928490490491u,1.5 5148.702890890891u,1.5 5148.703890890891u,0 5161.410911411411u,0 5161.411911411411u,1.5 5163.3659914914915u,1.5 5163.366991491492u,0 5164.343531531531u,0 5164.344531531531u,1.5 5173.1413918918915u,1.5 5173.142391891892u,0 5174.118931931932u,0 5174.119931931932u,1.5 5175.096471971972u,1.5 5175.0974719719725u,0 5181.939252252252u,0 5181.940252252252u,1.5 5182.9167922922925u,1.5 5182.917792292293u,0 5185.849412412412u,0 5185.850412412412u,1.5 5186.826952452452u,1.5 5186.827952452452u,0 5187.8044924924925u,0 5187.805492492493u,1.5 5197.5798928928925u,1.5 5197.580892892893u,0 5207.3552932932935u,0 5207.356293293294u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5209.310373373373u,0 5209.3113733733735u,1.5 5210.287913413413u,1.5 5210.288913413413u,0 5211.265453453453u,0 5211.266453453453u,1.5 5217.1306936936935u,1.5 5217.131693693694u,0 5218.108233733733u,0 5218.109233733733u,1.5 5219.085773773774u,1.5 5219.086773773774u,0 5220.063313813814u,0 5220.064313813814u,1.5 5221.040853853853u,1.5 5221.041853853853u,0 5228.861174174174u,0 5228.8621741741745u,1.5 5230.816254254254u,1.5 5230.817254254254u,0 5231.7937942942945u,0 5231.794794294295u,1.5 5239.614114614615u,1.5 5239.615114614615u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5257.209835335335u,1.5 5257.210835335335u,0 5258.187375375375u,0 5258.1883753753755u,1.5 5260.142455455456u,1.5 5260.143455455456u,0 5261.1199954954955u,0 5261.120995495496u,1.5 5262.097535535535u,1.5 5262.098535535535u,0 5264.052615615616u,0 5264.053615615616u,1.5 5265.030155655656u,1.5 5265.031155655656u,0 5271.872935935936u,0 5271.873935935936u,1.5 5274.805556056056u,1.5 5274.806556056056u,0 5275.783096096096u,0 5275.784096096097u,1.5 5281.648336336336u,1.5 5281.649336336336u,0 5282.625876376376u,0 5282.6268763763765u,1.5 5283.603416416417u,1.5 5283.604416416417u,0 5287.513576576576u,0 5287.5145765765765u,1.5 5288.491116616617u,1.5 5288.492116616617u,0 5292.401276776777u,0 5292.402276776777u,1.5 5303.154217217217u,1.5 5303.155217217217u,0 5313.907157657658u,0 5313.908157657658u,1.5 5315.862237737737u,1.5 5315.863237737737u,0 5316.839777777778u,0 5316.840777777778u,1.5 5327.592718218218u,1.5 5327.593718218218u,0 5339.323198698698u,0 5339.324198698699u,1.5 5346.165978978979u,1.5 5346.166978978979u,0 5347.143519019019u,0 5347.144519019019u,1.5 5349.098599099099u,1.5 5349.0995990991u,0 5350.076139139139u,0 5350.077139139139u,1.5 5352.031219219219u,1.5 5352.032219219219u,0 5359.851539539539u,0 5359.852539539539u,1.5 5360.829079579579u,1.5 5360.830079579579u,0 5365.71677977978u,0 5365.71777977978u,1.5 5376.46972022022u,1.5 5376.47072022022u,0 5377.447260260261u,0 5377.448260260261u,1.5 5378.4248003003u,1.5 5378.425800300301u,0 5380.37988038038u,0 5380.38088038038u,1.5 5381.357420420421u,1.5 5381.358420420421u,0 5392.110360860861u,0 5392.111360860861u,1.5 5393.0879009009u,1.5 5393.088900900901u,0 5396.020521021021u,0 5396.021521021021u,1.5 5411.661161661662u,1.5 5411.662161661662u,0 5412.638701701701u,0 5412.639701701702u,1.5 5415.571321821822u,1.5 5415.572321821822u,0 5417.526401901901u,0 5417.527401901902u,1.5 5418.503941941942u,1.5 5418.504941941942u,0 5433.167042542542u,0 5433.168042542542u,1.5 5434.144582582582u,1.5 5434.145582582582u,0 5435.122122622623u,0 5435.123122622623u,1.5 5436.099662662663u,1.5 5436.100662662663u,0 5437.077202702702u,0 5437.078202702703u,1.5 5442.942442942943u,1.5 5442.943442942943u,0 5443.919982982983u,0 5443.920982982983u,1.5 5457.605543543543u,1.5 5457.606543543543u,0 5458.583083583583u,0 5458.584083583583u,1.5 5460.538163663664u,1.5 5460.539163663664u,0 5461.515703703703u,0 5461.516703703704u,1.5 5466.403403903903u,1.5 5466.404403903904u,0 5467.380943943944u,0 5467.381943943944u,1.5 5468.358483983984u,1.5 5468.359483983984u,0 5469.336024024024u,0 5469.337024024024u,1.5 5471.291104104104u,1.5 5471.2921041041045u,0 5473.246184184184u,0 5473.247184184184u,1.5 5474.223724224224u,1.5 5474.224724224224u,0 5475.201264264265u,0 5475.202264264265u,1.5 5476.178804304304u,1.5 5476.1798043043045u,0 5478.133884384384u,0 5478.134884384384u,1.5 5479.1114244244245u,1.5 5479.112424424425u,0 5481.066504504504u,0 5481.0675045045045u,1.5 5482.044044544544u,1.5 5482.045044544544u,0 5490.841904904904u,0 5490.842904904905u,1.5 5491.819444944945u,1.5 5491.820444944945u,0 5493.774525025025u,0 5493.775525025025u,1.5 5494.752065065065u,1.5 5494.753065065065u,0 5497.684685185185u,0 5497.685685185185u,1.5 5498.662225225225u,1.5 5498.663225225225u,0 5511.370245745745u,0 5511.371245745745u,1.5 5512.347785785786u,1.5 5512.348785785786u,0 5520.168106106106u,0 5520.1691061061065u,1.5 5521.145646146146u,1.5 5521.146646146146u,0 5524.078266266267u,0 5524.079266266267u,1.5 5525.055806306306u,1.5 5525.0568063063065u,0 5527.9884264264265u,0 5527.989426426427u,1.5 5528.965966466467u,1.5 5528.966966466467u,0 5529.943506506506u,0 5529.9445065065065u,1.5 5533.853666666667u,1.5 5533.854666666667u,0 5534.831206706706u,0 5534.8322067067065u,1.5 5540.696446946947u,1.5 5540.697446946947u,0 5541.673986986987u,0 5541.674986986987u,1.5 5542.6515270270265u,1.5 5542.652527027027u,0 5543.629067067067u,0 5543.630067067067u,1.5 5557.3146276276275u,1.5 5557.315627627628u,0 5558.292167667668u,0 5558.293167667668u,1.5 5564.157407907907u,1.5 5564.1584079079075u,0 5568.067568068068u,0 5568.068568068068u,1.5 5569.045108108108u,1.5 5569.0461081081085u,0 5584.685748748749u,0 5584.686748748749u,1.5 5585.663288788789u,1.5 5585.664288788789u,0 5587.618368868869u,0 5587.619368868869u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5602.28146946947u,0 5602.28246946947u,1.5 5604.236549549549u,1.5 5604.237549549549u,0 5606.1916296296295u,0 5606.19262962963u,1.5 5607.16916966967u,1.5 5607.17016966967u,0 5616.94457007007u,0 5616.94557007007u,1.5 5617.92211011011u,1.5 5617.92311011011u,0 5619.87719019019u,0 5619.87819019019u,1.5 5620.8547302302295u,1.5 5620.85573023023u,0 5623.78735035035u,0 5623.78835035035u,1.5 5626.719970470471u,1.5 5626.720970470471u,0 5627.69751051051u,0 5627.6985105105105u,1.5 5637.47291091091u,1.5 5637.4739109109105u,0 5648.225851351351u,0 5648.226851351351u,1.5 5650.180931431431u,1.5 5650.181931431432u,0 5652.136011511511u,0 5652.137011511511u,1.5 5659.956331831831u,1.5 5659.957331831832u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5662.888951951952u,1.5 5662.889951951952u,0 5673.641892392392u,0 5673.642892392392u,1.5 5674.619432432432u,1.5 5674.620432432433u,0 5675.596972472473u,0 5675.597972472473u,1.5 5685.372372872873u,1.5 5685.373372872873u,0 5686.349912912912u,0 5686.3509129129125u,1.5 5687.327452952953u,1.5 5687.328452952953u,0 5696.125313313313u,0 5696.126313313313u,1.5 5698.080393393393u,1.5 5698.081393393393u,0 5699.057933433433u,0 5699.058933433434u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5719.586274274275u,0 5719.587274274275u,1.5 5728.384134634634u,1.5 5728.385134634635u,0 5729.361674674675u,0 5729.362674674675u,1.5 5730.339214714714u,1.5 5730.340214714714u,0 5739.137075075075u,0 5739.138075075075u,1.5 5740.114615115115u,1.5 5740.115615115115u,0 5741.092155155155u,0 5741.093155155155u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5760.6429559559565u,0 5760.643955955957u,1.5 5762.598036036035u,1.5 5762.599036036036u,0 5763.575576076076u,0 5763.576576076076u,1.5 5769.440816316316u,1.5 5769.441816316316u,0 5770.4183563563565u,0 5770.419356356357u,1.5 5771.395896396396u,1.5 5771.396896396396u,0 5780.1937567567575u,0 5780.194756756758u,1.5 5781.171296796797u,1.5 5781.172296796797u,0 5782.148836836836u,0 5782.149836836837u,1.5 5785.0814569569575u,1.5 5785.082456956958u,0 5786.058996996997u,0 5786.059996996997u,1.5 5791.924237237236u,1.5 5791.925237237237u,0 5794.8568573573575u,0 5794.857857357358u,1.5 5795.834397397397u,1.5 5795.835397397397u,0 5802.677177677678u,0 5802.678177677678u,1.5 5803.654717717717u,1.5 5803.655717717717u,0 5804.632257757758u,0 5804.633257757759u,1.5 5811.475038038037u,1.5 5811.476038038038u,0 5812.452578078078u,0 5812.453578078078u,1.5 5814.4076581581585u,1.5 5814.408658158159u,0 5816.362738238237u,0 5816.363738238238u,1.5 5817.340278278279u,1.5 5817.341278278279u,0 5827.115678678679u,0 5827.116678678679u,1.5 5833.958458958959u,1.5 5833.95945895896u,0 5834.935998998999u,0 5834.936998998999u,1.5 5836.891079079079u,1.5 5836.892079079079u,0 5837.868619119119u,0 5837.869619119119u,1.5 5839.823699199199u,1.5 5839.824699199199u,0 5849.5990995996u,0 5849.6000995996u,1.5 5850.576639639639u,1.5 5850.5776396396395u,0 5851.55417967968u,0 5851.55517967968u,1.5 5861.32958008008u,1.5 5861.33058008008u,0 5862.30712012012u,0 5862.30812012012u,1.5 5863.2846601601605u,1.5 5863.285660160161u,0 5864.2622002002u,0 5864.2632002002u,1.5 5865.239740240239u,1.5 5865.24074024024u,0 5866.217280280281u,0 5866.218280280281u,1.5 5867.19482032032u,1.5 5867.19582032032u,0 5877.947760760761u,0 5877.948760760762u,1.5 5878.925300800801u,1.5 5878.926300800801u,0 5879.90284084084u,0 5879.9038408408405u,1.5 5880.880380880881u,1.5 5880.881380880881u,0 5881.857920920921u,0 5881.858920920921u,1.5 5891.633321321321u,1.5 5891.634321321321u,0 5892.6108613613615u,0 5892.611861361362u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5896.521021521521u,0 5896.522021521521u,1.5 5897.4985615615615u,1.5 5897.499561561562u,0 5907.273961961962u,0 5907.274961961963u,1.5 5908.251502002002u,1.5 5908.252502002002u,0 5910.206582082082u,0 5910.207582082082u,1.5 5911.184122122122u,1.5 5911.185122122122u,0 5913.139202202202u,0 5913.140202202202u,1.5 5930.734922922923u,1.5 5930.735922922923u,0 5931.712462962963u,0 5931.713462962964u,1.5 5935.622623123123u,1.5 5935.623623123123u,0 5942.465403403403u,0 5942.466403403403u,1.5 5943.442943443443u,1.5 5943.4439434434435u,0 5962.993744244243u,0 5962.9947442442435u,1.5 5963.971284284285u,1.5 5963.972284284285u,0 5964.948824324324u,0 5964.949824324324u,1.5 5965.926364364364u,1.5 5965.927364364365u,0 5967.881444444444u,0 5967.882444444444u,1.5 5968.858984484485u,1.5 5968.859984484485u,0 5970.814064564564u,0 5970.815064564565u,1.5 5971.791604604605u,1.5 5971.792604604605u,0 5972.769144644644u,0 5972.7701446446445u,1.5 5973.746684684685u,1.5 5973.747684684685u,0 5974.724224724724u,0 5974.725224724724u,1.5 5976.679304804805u,1.5 5976.680304804805u,0 5977.656844844844u,0 5977.6578448448445u,1.5 5980.589464964965u,1.5 5980.590464964966u,0 5981.567005005005u,0 5981.568005005005u,1.5 5994.275025525525u,1.5 5994.276025525525u,0 5995.252565565565u,0 5995.253565565566u,1.5 6001.117805805806u,1.5 6001.118805805806u,0 6002.095345845845u,0 6002.0963458458455u,1.5 6013.825826326326u,1.5 6013.826826326326u,0 6014.803366366366u,0 6014.804366366367u,1.5 6019.691066566566u,1.5 6019.692066566567u,0 6020.668606606607u,0 6020.669606606607u,1.5 6024.578766766767u,1.5 6024.5797667667675u,0 6025.556306806807u,0 6025.557306806807u,1.5 6029.466466966967u,1.5 6029.467466966968u,0 6031.421547047046u,0 6031.4225470470465u,1.5 6033.376627127127u,1.5 6033.377627127127u,0 6034.354167167167u,0 6034.355167167168u,1.5 6035.331707207207u,1.5 6035.332707207207u,0 6037.286787287288u,0 6037.287787287288u,1.5 6038.264327327327u,1.5 6038.265327327327u,0 6061.7252882882885u,0 6061.726288288289u,1.5 6063.680368368368u,1.5 6063.681368368369u,0 6064.657908408408u,0 6064.658908408408u,1.5 6065.635448448448u,1.5 6065.636448448448u,0 6066.612988488489u,0 6066.613988488489u,1.5 6074.433308808809u,1.5 6074.434308808809u,0 6075.410848848848u,0 6075.411848848848u,1.5 6082.253629129129u,1.5 6082.254629129129u,0 6083.231169169169u,0 6083.2321691691695u,1.5 6084.208709209209u,1.5 6084.209709209209u,0 6085.186249249249u,0 6085.187249249249u,1.5 6087.141329329329u,1.5 6087.142329329329u,0 6088.118869369369u,0 6088.11986936937u,1.5 6090.073949449449u,1.5 6090.074949449449u,0 6091.0514894894895u,0 6091.05248948949u,1.5 6092.029029529529u,1.5 6092.030029529529u,0 6103.75951001001u,0 6103.76051001001u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6120.3776906906905u,1.5 6120.378690690691u,0 6121.35523073073u,0 6121.35623073073u,1.5 6122.332770770771u,1.5 6122.3337707707715u,0 6123.310310810811u,0 6123.311310810811u,1.5 6124.28785085085u,1.5 6124.28885085085u,0 6133.085711211211u,0 6133.086711211211u,1.5 6134.063251251251u,1.5 6134.064251251251u,0 6136.995871371371u,0 6136.9968713713715u,1.5 6147.748811811812u,1.5 6147.749811811812u,0 6148.726351851851u,0 6148.727351851851u,1.5 6149.7038918918915u,1.5 6149.704891891892u,0 6151.658971971972u,0 6151.6599719719725u,1.5 6152.636512012012u,1.5 6152.637512012012u,0 6160.456832332332u,0 6160.457832332332u,1.5 6161.434372372372u,1.5 6161.4353723723725u,0 6162.411912412412u,0 6162.412912412412u,1.5 6163.389452452452u,1.5 6163.390452452452u,0 6164.3669924924925u,0 6164.367992492493u,1.5 6172.187312812813u,1.5 6172.188312812813u,0 6173.164852852852u,0 6173.165852852852u,1.5 6175.119932932933u,1.5 6175.120932932933u,0 6186.850413413413u,0 6186.851413413413u,1.5 6195.648273773774u,1.5 6195.649273773774u,0 6196.625813813814u,0 6196.626813813814u,1.5 6197.603353853853u,1.5 6197.604353853853u,0 6207.378754254254u,0 6207.379754254254u,1.5 6217.154154654654u,1.5 6217.155154654654u,0 6219.109234734734u,0 6219.110234734734u,1.5 6220.086774774775u,1.5 6220.087774774775u,0 6229.862175175175u,0 6229.8631751751755u,1.5 6230.839715215215u,1.5 6230.840715215215u,0 6231.817255255255u,0 6231.818255255255u,1.5 6238.660035535535u,1.5 6238.661035535535u,0 6239.637575575575u,0 6239.6385755755755u,1.5 6240.615115615616u,1.5 6240.616115615616u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6251.368056056055u,1.5 6251.369056056055u,0 6252.345596096096u,0 6252.346596096097u,1.5 6259.188376376376u,1.5 6259.1893763763765u,0 6260.165916416417u,0 6260.166916416417u,1.5 6261.143456456457u,1.5 6261.144456456457u,0 6262.120996496496u,0 6262.121996496497u,1.5 6263.098536536536u,1.5 6263.099536536536u,0 6267.0086966966965u,0 6267.009696696697u,1.5 6267.986236736736u,1.5 6267.987236736736u,0 6271.8963968968965u,0 6271.897396896897u,1.5 6279.716717217217u,1.5 6279.717717217217u,0 6280.694257257258u,0 6280.695257257258u,1.5 6281.671797297297u,1.5 6281.672797297298u,0 6282.649337337337u,0 6282.650337337337u,1.5 6283.626877377377u,1.5 6283.627877377377u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6293.402277777778u,0 6293.403277777778u,1.5 6303.177678178178u,1.5 6303.178678178178u,0 6315.885698698698u,0 6315.886698698699u,1.5 6323.706019019019u,1.5 6323.707019019019u,0 6324.683559059059u,0 6324.684559059059u,1.5 6325.661099099099u,1.5 6325.6620990991u,0 6326.638639139139u,0 6326.639639139139u,1.5 6327.616179179179u,1.5 6327.617179179179u,0 6338.36911961962u,0 6338.37011961962u,1.5 6350.0996001001u,1.5 6350.100600100101u,0 6351.07714014014u,0 6351.07814014014u,1.5 6352.05468018018u,1.5 6352.05568018018u,0 6355.96484034034u,0 6355.96584034034u,1.5 6356.94238038038u,1.5 6356.94338038038u,0 6361.83008058058u,0 6361.83108058058u,1.5 6362.807620620621u,1.5 6362.808620620621u,0 6364.7627007007u,0 6364.763700700701u,1.5 6367.695320820821u,1.5 6367.696320820821u,0 6368.672860860861u,0 6368.673860860861u,1.5 6375.515641141141u,1.5 6375.516641141141u,0 6376.493181181181u,0 6376.494181181181u,1.5 6378.448261261262u,1.5 6378.449261261262u,0 6381.380881381381u,0 6381.381881381381u,1.5 6382.358421421422u,1.5 6382.359421421422u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6393.111361861862u,0 6393.112361861862u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6396.043981981982u,1.5 6396.044981981982u,0 6397.021522022022u,0 6397.022522022022u,1.5 6411.684622622623u,1.5 6411.685622622623u,0 6412.662162662663u,0 6412.663162662663u,1.5 6413.639702702702u,1.5 6413.640702702703u,0 6414.617242742742u,0 6414.618242742742u,1.5 6416.572322822823u,1.5 6416.573322822823u,0 6420.482482982983u,0 6420.483482982983u,1.5 6421.460023023023u,1.5 6421.461023023023u,0 6427.325263263264u,0 6427.326263263264u,1.5 6428.302803303303u,1.5 6428.3038033033035u,0 6432.212963463464u,0 6432.213963463464u,1.5 6433.190503503503u,1.5 6433.191503503504u,0 6434.168043543543u,0 6434.169043543543u,1.5 6435.145583583583u,1.5 6435.146583583583u,0 6436.1231236236235u,0 6436.124123623624u,1.5 6438.078203703703u,1.5 6438.079203703704u,0 6439.055743743743u,0 6439.056743743743u,1.5 6442.965903903903u,1.5 6442.966903903904u,0 6443.943443943944u,0 6443.944443943944u,1.5 6460.5616246246245u,1.5 6460.562624624625u,0 6461.539164664665u,0 6461.540164664665u,1.5 6466.426864864865u,1.5 6466.427864864865u,0 6467.404404904904u,0 6467.405404904905u,1.5 6468.381944944945u,1.5 6468.382944944945u,0 6469.359484984985u,0 6469.360484984985u,1.5 6470.337025025025u,1.5 6470.338025025025u,0 6471.314565065065u,0 6471.315565065065u,1.5 6472.292105105105u,1.5 6472.2931051051055u,0 6473.269645145145u,0 6473.270645145145u,1.5 6474.247185185185u,1.5 6474.248185185185u,0 6477.179805305305u,0 6477.1808053053055u,1.5 6478.157345345345u,1.5 6478.158345345345u,0 6483.045045545545u,0 6483.046045545545u,1.5 6484.022585585586u,1.5 6484.023585585586u,0 6485.0001256256255u,0 6485.001125625626u,1.5 6485.977665665666u,1.5 6485.978665665666u,0 6486.955205705705u,0 6486.9562057057055u,1.5 6487.932745745745u,1.5 6487.933745745745u,0 6489.8878258258255u,0 6489.888825825826u,1.5 6490.865365865866u,1.5 6490.866365865866u,0 6494.775526026026u,0 6494.776526026026u,1.5 6495.753066066066u,1.5 6495.754066066066u,0 6502.595846346346u,0 6502.596846346346u,1.5 6503.573386386386u,1.5 6503.574386386386u,0 6504.5509264264265u,0 6504.551926426427u,1.5 6505.528466466467u,1.5 6505.529466466467u,0 6509.4386266266265u,0 6509.439626626627u,1.5 6510.416166666667u,1.5 6510.417166666667u,0 6512.371246746747u,0 6512.372246746747u,1.5 6513.348786786787u,1.5 6513.349786786787u,0 6514.3263268268265u,0 6514.327326826827u,1.5 6515.303866866867u,1.5 6515.304866866867u,0 6516.281406906906u,0 6516.2824069069065u,1.5 6517.258946946947u,1.5 6517.259946946947u,0 6519.2140270270265u,0 6519.215027027027u,1.5 6520.191567067067u,1.5 6520.192567067067u,0 6521.169107107107u,0 6521.1701071071075u,1.5 6522.146647147147u,1.5 6522.147647147147u,0 6523.124187187187u,0 6523.125187187187u,1.5 6524.101727227227u,1.5 6524.102727227227u,0 6525.079267267268u,0 6525.080267267268u,1.5 6526.056807307307u,1.5 6526.0578073073075u,0 6528.011887387387u,0 6528.012887387387u,1.5 6529.966967467468u,1.5 6529.967967467468u,0 6531.922047547547u,0 6531.923047547547u,1.5 6532.899587587588u,1.5 6532.900587587588u,0 6533.8771276276275u,0 6533.878127627628u,1.5 6534.854667667668u,1.5 6534.855667667668u,0 6535.832207707707u,0 6535.8332077077075u,1.5 6538.7648278278275u,1.5 6538.765827827828u,0 6539.742367867868u,0 6539.743367867868u,1.5 6557.338088588589u,1.5 6557.339088588589u,0 6558.3156286286285u,0 6558.316628628629u,1.5 6560.270708708708u,1.5 6560.2717087087085u,0 6561.248248748749u,0 6561.249248748749u,1.5 6562.225788788789u,1.5 6562.226788788789u,0 6563.2033288288285u,0 6563.204328828829u,1.5 6564.180868868869u,1.5 6564.181868868869u,0 6566.135948948949u,0 6566.136948948949u,1.5 6567.113488988989u,1.5 6567.114488988989u,0 6571.023649149149u,0 6571.024649149149u,1.5 6572.001189189189u,1.5 6572.002189189189u,0 6584.709209709709u,0 6584.7102097097095u,1.5 6585.68674974975u,1.5 6585.68774974975u,0 6586.66428978979u,0 6586.66528978979u,1.5 6588.61936986987u,1.5 6588.62036986987u,0 6591.55198998999u,0 6591.55298998999u,1.5 6602.30493043043u,1.5 6602.305930430431u,0 6603.282470470471u,0 6603.283470470471u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6608.170170670671u,0 6608.171170670671u,1.5 6609.14771071071u,1.5 6609.1487107107105u,0 6619.900651151151u,0 6619.901651151151u,1.5 6620.878191191191u,1.5 6620.879191191191u,0 6622.833271271272u,0 6622.834271271272u,1.5 6623.810811311311u,1.5 6623.811811311311u,0 6624.788351351351u,0 6624.789351351351u,1.5 6632.608671671672u,1.5 6632.609671671672u,0 6633.586211711711u,0 6633.5872117117115u,1.5 6634.563751751752u,1.5 6634.564751751752u,0 6635.541291791792u,0 6635.542291791792u,1.5 6636.518831831831u,1.5 6636.519831831832u,0 6640.428991991992u,0 6640.429991991992u,1.5 6641.4065320320315u,1.5 6641.407532032032u,0 6650.204392392392u,0 6650.205392392392u,1.5 6652.159472472473u,1.5 6652.160472472473u,0 6653.137012512512u,0 6653.138012512512u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6671.710273273274u,0 6671.711273273274u,1.5 6672.687813313313u,1.5 6672.688813313313u,0 6674.642893393393u,0 6674.643893393393u,1.5 6676.597973473474u,1.5 6676.598973473474u,0 6677.575513513513u,0 6677.576513513513u,1.5 6684.418293793794u,1.5 6684.419293793794u,0 6685.395833833833u,0 6685.396833833834u,1.5 6687.350913913913u,1.5 6687.351913913913u,0 6697.126314314314u,0 6697.127314314314u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6716.677115115115u,0 6716.678115115115u,1.5 6717.654655155155u,1.5 6717.655655155155u,0 6719.609735235234u,0 6719.610735235235u,1.5 6720.587275275276u,1.5 6720.588275275276u,0 6721.564815315315u,0 6721.565815315315u,1.5 6722.542355355355u,1.5 6722.543355355355u,0 6723.519895395395u,0 6723.520895395395u,1.5 6725.474975475476u,1.5 6725.475975475476u,0 6726.452515515515u,0 6726.453515515515u,1.5 6729.385135635635u,1.5 6729.386135635636u,0 6730.362675675676u,0 6730.363675675676u,1.5 6731.340215715715u,1.5 6731.341215715715u,0 6739.160536036035u,0 6739.161536036036u,1.5 6740.138076076076u,1.5 6740.139076076076u,0 6741.115616116116u,0 6741.116616116116u,1.5 6747.958396396396u,1.5 6747.959396396396u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6756.7562567567575u,0 6756.757256756758u,1.5 6757.733796796797u,1.5 6757.734796796797u,0 6758.711336836836u,0 6758.712336836837u,1.5 6759.688876876877u,1.5 6759.689876876877u,0 6762.621496996997u,0 6762.622496996997u,1.5 6770.441817317317u,1.5 6770.442817317317u,0 6772.396897397397u,0 6772.397897397397u,1.5 6773.374437437437u,1.5 6773.3754374374375u,0 6780.217217717717u,0 6780.218217717717u,1.5 6792.925238238237u,1.5 6792.926238238238u,0 6802.700638638638u,0 6802.7016386386385u,1.5 6804.655718718718u,1.5 6804.656718718718u,0 6805.633258758759u,0 6805.63425875876u,1.5 6812.476039039038u,1.5 6812.477039039039u,0 6813.453579079079u,0 6813.454579079079u,1.5 6816.386199199199u,1.5 6816.387199199199u,0 6824.206519519519u,0 6824.207519519519u,1.5 6825.1840595595595u,1.5 6825.18505955956u,0 6826.1615995996u,0 6826.1625995996u,1.5 6827.139139639639u,1.5 6827.1401396396395u,0 6828.11667967968u,0 6828.11767967968u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6846.68994044044u,0 6846.6909404404405u,1.5 6847.667480480481u,1.5 6847.668480480481u,0 6850.600100600601u,0 6850.601100600601u,1.5 6854.510260760761u,1.5 6854.511260760762u,0 6855.487800800801u,0 6855.488800800801u,1.5 6864.285661161161u,1.5 6864.286661161162u,0 6865.263201201201u,0 6865.264201201201u,1.5 6866.24074124124u,1.5 6866.241741241241u,0 6873.083521521521u,0 6873.084521521521u,1.5 6874.0610615615615u,1.5 6874.062061561562u,0 6877.971221721721u,0 6877.972221721721u,1.5 6878.948761761762u,1.5 6878.949761761763u,0 6879.926301801802u,0 6879.927301801802u,1.5 6891.656782282283u,1.5 6891.657782282283u,0 6892.634322322322u,0 6892.635322322322u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6911.207583083083u,0 6911.208583083083u,1.5 6912.185123123123u,1.5 6912.186123123123u,0 6913.162663163163u,0 6913.163663163164u,1.5 6915.117743243242u,1.5 6915.1187432432425u,0 6916.095283283284u,0 6916.096283283284u,1.5 6929.780843843843u,1.5 6929.7818438438435u,0 6930.758383883884u,0 6930.759383883884u,1.5 6935.646084084084u,1.5 6935.647084084084u,0 6937.601164164164u,0 6937.602164164165u,1.5 6938.578704204204u,1.5 6938.579704204204u,0 6943.466404404404u,0 6943.467404404404u,1.5 6944.443944444444u,1.5 6944.444944444444u,0 6957.151964964965u,0 6957.152964964966u,1.5 6958.129505005005u,1.5 6958.130505005005u,0 6963.994745245244u,0 6963.9957452452445u,1.5 6964.972285285286u,1.5 6964.973285285286u,0 6965.949825325325u,0 6965.950825325325u,1.5 6966.927365365365u,1.5 6966.928365365366u,0 6968.882445445445u,0 6968.883445445445u,1.5 6971.815065565565u,1.5 6971.816065565566u,0 6972.792605605606u,0 6972.793605605606u,1.5 6973.770145645645u,1.5 6973.771145645645u,0 6974.747685685686u,0 6974.748685685686u,1.5 6975.725225725725u,1.5 6975.726225725725u,0 6976.702765765766u,0 6976.703765765767u,1.5 6980.612925925926u,1.5 6980.613925925926u,0 6981.590465965966u,0 6981.591465965967u,1.5 6986.478166166166u,1.5 6986.479166166167u,0 6987.455706206206u,0 6987.456706206206u,1.5 6988.433246246245u,1.5 6988.4342462462455u,0 6989.410786286287u,0 6989.411786286287u,1.5 6990.388326326326u,1.5 6990.389326326326u,0 6991.365866366366u,0 6991.366866366367u,1.5
vbb23 bb23 0 pwl 0,1.5  61.58452252252251u,1.5 61.58552252252252u,0 62.56206256256256u,0 62.563062562562564u,1.5 63.539602602602606u,1.5 63.54060260260261u,0 64.51714264264264u,0 64.51814264264264u,1.5 65.49468268268268u,1.5 65.49568268268268u,0 66.47222272272272u,0 66.47322272272272u,1.5 67.44976276276276u,1.5 67.45076276276276u,0 68.4273028028028u,0 68.4283028028028u,1.5 69.40484284284284u,1.5 69.40584284284284u,0 70.38238288288288u,0 70.38338288288288u,1.5 71.35992292292292u,1.5 71.36092292292292u,0 107.5289044044044u,0 107.5299044044044u,1.5 134.90002552552554u,1.5 134.9010255255255u,0 135.8775655655656u,0 135.87856556556557u,1.5 137.83264564564567u,1.5 137.83364564564565u,0 163.2486866866867u,0 163.2496866866867u,1.5 184.7545675675676u,1.5 184.75556756756757u,0 186.70964764764764u,0 186.71064764764762u,1.5 187.6871876876877u,1.5 187.68818768768767u,0 208.21552852852852u,0 208.2165285285285u,1.5 225.81124924924927u,1.5 225.81224924924925u,0 226.7887892892893u,0 226.78978928928927u,1.5 228.74386936936938u,1.5 228.74486936936935u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 271.75563113113117u,1.5 271.75663113113114u,0 291.3064319319319u,0 291.3074319319319u,1.5 292.28397197197194u,1.5 292.2849719719719u,0 294.23905205205205u,0 294.240052052052u,1.5 314.76739289289293u,1.5 314.7683928928929u,0 316.722472972973u,0 316.72347297297296u,1.5 317.700013013013u,1.5 317.701013013013u,0 334.31819369369373u,0 334.3191936936937u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 337.2508138138138u,0 337.2518138138138u,1.5 362.6668548548549u,1.5 362.66785485485485u,0 363.6443948948949u,0 363.6453948948949u,1.5 364.621934934935u,1.5 364.62293493493496u,0 391.99305605605605u,0 391.994056056056u,1.5 392.9705960960961u,1.5 392.97159609609605u,0 394.9256761761762u,0 394.92667617617616u,1.5 396.8807562562563u,1.5 396.88175625625627u,0 397.85829629629626u,0 397.85929629629624u,1.5 434.0272777777778u,1.5 434.02827777777776u,0 435.98235785785783u,0 435.9833578578578u,1.5 436.9598978978979u,1.5 436.9608978978979u,0 442.82513813813813u,0 442.8261381381381u,1.5 443.80267817817816u,1.5 443.80367817817813u,0 447.7128383383383u,0 447.7138383383383u,1.5 448.69037837837834u,1.5 448.6913783783783u,0 560.1299429429429u,0 560.1309429429429u,1.5 562.085023023023u,1.5 562.086023023023u,0 565.0176431431431u,0 565.0186431431431u,1.5 565.9951831831833u,1.5 565.9961831831832u,0 566.9727232232233u,0 566.9737232232233u,1.5 567.9502632632633u,1.5 567.9512632632633u,0 568.9278033033033u,0 568.9288033033033u,1.5 605.0967847847849u,1.5 605.0977847847848u,0 607.0518648648649u,0 607.0528648648649u,1.5 608.0294049049048u,1.5 608.0304049049048u,0 633.445445945946u,0 633.4464459459459u,1.5 634.422985985986u,1.5 634.423985985986u,0 635.400526026026u,0 635.401526026026u,1.5 636.378066066066u,1.5 636.379066066066u,0 637.355606106106u,0 637.356606106106u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 664.7267272272272u,0 664.7277272272272u,1.5 665.7042672672673u,1.5 665.7052672672672u,0 684.277528028028u,0 684.278528028028u,1.5 687.2101481481482u,1.5 687.2111481481481u,0 688.1876881881882u,0 688.1886881881882u,1.5 704.8058688688689u,1.5 704.8068688688688u,0 705.783408908909u,0 705.784408908909u,1.5 708.716029029029u,1.5 708.7170290290289u,0 727.2892897897898u,0 727.2902897897898u,1.5 728.2668298298298u,1.5 728.2678298298298u,0 730.22190990991u,0 730.22290990991u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 770.3010515515515u,0 770.3020515515515u,1.5 791.8069324324325u,1.5 791.8079324324325u,0 813.3128133133133u,0 813.3138133133133u,1.5 815.2678933933934u,1.5 815.2688933933933u,0 816.2454334334335u,0 816.2464334334335u,1.5 817.2229734734735u,1.5 817.2239734734735u,0 818.2005135135136u,0 818.2015135135135u,1.5 834.8186941941941u,1.5 834.8196941941941u,0 835.7962342342342u,0 835.7972342342342u,1.5 836.7737742742743u,1.5 836.7747742742743u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 861.2122752752753u,0 861.2132752752752u,1.5 862.1898153153153u,1.5 862.1908153153153u,0 863.1673553553553u,0 863.1683553553553u,1.5 865.1224354354355u,1.5 865.1234354354355u,0 866.0999754754755u,0 866.1009754754755u,1.5 895.4261766766766u,1.5 895.4271766766766u,0 929.6400780780781u,0 929.6410780780781u,1.5 930.6176181181181u,1.5 930.6186181181181u,0 934.5277782782782u,0 934.5287782782782u,1.5 935.5053183183182u,1.5 935.5063183183182u,0 936.4828583583584u,0 936.4838583583584u,1.5 939.4154784784785u,1.5 939.4164784784784u,0 940.3930185185185u,0 940.3940185185185u,1.5 1063.5630635635634u,1.5 1063.5640635635636u,0 1066.4956836836834u,0 1066.4966836836836u,1.5 1067.4732237237235u,1.5 1067.4742237237238u,0 1106.5748253253253u,0 1106.5758253253255u,1.5 1135.9010265265265u,1.5 1135.9020265265267u,0 1136.8785665665666u,0 1136.8795665665668u,1.5 1137.8561066066065u,1.5 1137.8571066066067u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1182.8229484484484u,1.5 1182.8239484484486u,0 1183.8004884884883u,0 1183.8014884884885u,1.5 1184.7780285285285u,1.5 1184.7790285285287u,0 1185.7555685685686u,0 1185.7565685685688u,1.5 1186.7331086086085u,1.5 1186.7341086086087u,0 1207.2614494494494u,0 1207.2624494494496u,1.5 1227.7897902902903u,1.5 1227.7907902902905u,0 1229.7448703703703u,0 1229.7458703703705u,1.5 1230.7224104104102u,1.5 1230.7234104104105u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1268.8464719719718u,1.5 1268.847471971972u,0 1269.8240120120117u,0 1269.825012012012u,1.5 1272.756632132132u,1.5 1272.7576321321321u,0 1289.3748128128127u,0 1289.375812812813u,1.5 1290.3523528528526u,1.5 1290.3533528528528u,0 1293.2849729729728u,0 1293.285972972973u,1.5 1294.2625130130127u,1.5 1294.263513013013u,0 1295.2400530530529u,0 1295.241053053053u,1.5 1314.7908538538536u,1.5 1314.7918538538538u,0 1336.2967347347346u,0 1336.2977347347348u,1.5 1337.2742747747748u,1.5 1337.275274774775u,0 1338.251814814815u,0 1338.252814814815u,1.5 1340.2068948948947u,1.5 1340.207894894895u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1361.7127757757758u,1.5 1361.713775775776u,0 1362.690315815816u,0 1362.691315815816u,1.5 1363.6678558558558u,1.5 1363.668855855856u,0 1364.6453958958957u,0 1364.646395895896u,1.5 1365.6229359359356u,1.5 1365.6239359359358u,0 1391.0389769769768u,0 1391.039976976977u,1.5 1392.016517017017u,1.5 1392.017517017017u,0 1392.9940570570568u,0 1392.995057057057u,1.5 1393.971597097097u,1.5 1393.9725970970972u,0 1394.9491371371369u,0 1394.950137137137u,1.5 1395.926677177177u,1.5 1395.9276771771772u,0 1396.9042172172171u,0 1396.9052172172173u,1.5 1436.9833588588588u,1.5 1436.984358858859u,0 1439.915978978979u,0 1439.9169789789792u,1.5 1440.8935190190189u,1.5 1440.894519019019u,0 1441.8710590590588u,0 1441.872059059059u,1.5 1442.848599099099u,1.5 1442.8495990990991u,0 1448.7138393393393u,0 1448.7148393393395u,1.5 1449.6913793793792u,1.5 1449.6923793793794u,0 1561.130943943944u,0 1561.1319439439442u,1.5 1562.108483983984u,1.5 1562.109483983984u,0 1564.063564064064u,0 1564.0645640640641u,1.5 1566.018644144144u,1.5 1566.0196441441442u,0 1566.996184184184u,0 1566.997184184184u,1.5 1601.2100855855854u,1.5 1601.2110855855856u,0 1602.1876256256255u,0 1602.1886256256257u,1.5 1605.1202457457457u,1.5 1605.121245745746u,0 1606.0977857857856u,0 1606.0987857857858u,1.5 1608.052865865866u,1.5 1608.053865865866u,0 1609.0304059059058u,0 1609.031405905906u,1.5 1610.007945945946u,1.5 1610.0089459459462u,0 1633.4689069069068u,0 1633.469906906907u,1.5 1634.446446946947u,1.5 1634.4474469469471u,0 1636.401527027027u,0 1636.4025270270272u,1.5 1637.3790670670671u,1.5 1637.3800670670673u,0 1638.356607107107u,0 1638.3576071071072u,1.5 1639.3341471471472u,1.5 1639.3351471471474u,0 1640.311687187187u,0 1640.3126871871873u,1.5 1658.884947947948u,1.5 1658.8859479479481u,0 1659.8624879879878u,0 1659.863487987988u,1.5 1663.7726481481482u,1.5 1663.7736481481484u,0 1685.278529029029u,0 1685.2795290290292u,1.5 1686.256069069069u,1.5 1686.2570690690693u,0 1687.233609109109u,0 1687.2346091091092u,1.5 1706.7844099099098u,1.5 1706.78540990991u,0 1707.76194994995u,0 1707.76294994995u,1.5 1708.73948998999u,1.5 1708.7404899899902u,0 1711.67211011011u,0 1711.6731101101102u,1.5 1712.6496501501501u,1.5 1712.6506501501503u,0 1725.3576706706706u,0 1725.3586706706708u,1.5 1726.3352107107105u,1.5 1726.3362107107107u,0 1730.2453708708708u,0 1730.246370870871u,1.5 1731.2229109109107u,1.5 1731.223910910911u,0 1732.2004509509509u,0 1732.201450950951u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1770.3245125125122u,0 1770.3255125125124u,1.5 1772.2795925925925u,1.5 1772.2805925925927u,0 1773.2571326326324u,0 1773.2581326326326u,1.5 1774.2346726726726u,1.5 1774.2356726726728u,0 1775.2122127127125u,0 1775.2132127127127u,1.5 1791.8303933933933u,1.5 1791.8313933933935u,0 1792.8079334334332u,0 1792.8089334334334u,1.5 1793.7854734734733u,1.5 1793.7864734734735u,0 1811.3811941941942u,0 1811.3821941941944u,1.5 1812.3587342342341u,1.5 1812.3597342342343u,0 1813.3362742742743u,0 1813.3372742742745u,1.5 1814.3138143143142u,1.5 1814.3148143143144u,0 1815.2913543543543u,0 1815.2923543543545u,1.5 1834.842155155155u,1.5 1834.8431551551553u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1861.235736236236u,0 1861.2367362362363u,1.5 1862.2132762762762u,1.5 1862.2142762762765u,0 1865.1458963963964u,0 1865.1468963963966u,1.5 1887.6293173173174u,1.5 1887.6303173173176u,0 1888.6068573573573u,0 1888.6078573573575u,1.5 1890.5619374374373u,1.5 1890.5629374374375u,0 1891.5394774774772u,0 1891.5404774774775u,1.5 1893.4945575575573u,1.5 1893.4955575575575u,0 1894.4720975975974u,0 1894.4730975975976u,1.5 1895.4496376376374u,1.5 1895.4506376376376u,0 1931.618619119119u,0 1931.6196191191193u,1.5 1932.596159159159u,1.5 1932.5971591591592u,0 1934.551239239239u,0 1934.5522392392393u,1.5 1936.5063193193193u,1.5 1936.5073193193195u,0 1937.4838593593593u,0 1937.4848593593595u,1.5 1938.4613993993994u,1.5 1938.4623993993996u,0 1939.4389394394395u,0 1939.4399394394397u,1.5 2058.698824324324u,1.5 2058.6998243243243u,0 2059.676364364364u,0 2059.677364364364u,1.5 2061.6314444444442u,1.5 2061.6324444444444u,0 2062.6089844844846u,0 2062.609984484485u,1.5 2064.5640645645644u,1.5 2064.5650645645646u,0 2065.5416046046043u,0 2065.5426046046045u,1.5 2066.5191446446447u,1.5 2066.520144644645u,0 2068.4742247247245u,0 2068.4752247247247u,1.5 2069.4517647647644u,1.5 2069.4527647647647u,0 2072.384384884885u,0 2072.3853848848853u,1.5 2073.3619249249246u,1.5 2073.3629249249248u,0 2104.643206206206u,0 2104.644206206206u,1.5 2107.575826326326u,1.5 2107.576826326326u,0 2108.553366366366u,0 2108.554366366366u,1.5 2112.463526526526u,1.5 2112.4645265265262u,0 2113.4410665665664u,0 2113.4420665665666u,1.5 2136.9020275275275u,1.5 2136.9030275275277u,0 2161.3405285285285u,0 2161.3415285285287u,1.5 2166.228228728729u,1.5 2166.229228728729u,0 2167.2057687687684u,0 2167.2067687687686u,1.5 2186.7565695695694u,1.5 2186.7575695695696u,0 2206.30737037037u,0 2206.30837037037u,1.5 2207.2849104104102u,1.5 2207.2859104104105u,0 2209.2399904904905u,0 2209.2409904904907u,1.5 2229.7683313313314u,1.5 2229.7693313313316u,0 2232.700951451451u,0 2232.7019514514514u,1.5 2233.6784914914915u,1.5 2233.6794914914917u,0 2250.296672172172u,0 2250.297672172172u,1.5 2270.8250130130127u,1.5 2270.826013013013u,0 2271.802553053053u,0 2271.8035530530533u,1.5 2272.780093093093u,1.5 2272.781093093093u,0 2291.3533538538536u,0 2291.354353853854u,1.5 2292.330893893894u,1.5 2292.331893893894u,0 2294.285973973974u,0 2294.286973973974u,1.5 2313.8367747747743u,1.5 2313.8377747747745u,0 2317.746934934935u,0 2317.747934934935u,1.5 2318.724474974975u,1.5 2318.725474974975u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2360.7586966966965u,1.5 2360.7596966966967u,0 2361.736236736737u,0 2361.737236736737u,1.5 2363.6913168168167u,1.5 2363.692316816817u,0 2364.6688568568566u,0 2364.6698568568568u,1.5 2365.646396896897u,1.5 2365.647396896897u,0 2388.1298178178176u,0 2388.130817817818u,1.5 2389.1073578578576u,1.5 2389.1083578578578u,0 2393.0175180180177u,0 2393.018518018018u,1.5 2393.995058058058u,1.5 2393.996058058058u,0 2394.972598098098u,0 2394.973598098098u,1.5 2395.9501381381383u,1.5 2395.9511381381385u,0 2396.927678178178u,0 2396.9286781781784u,1.5 2398.882758258258u,1.5 2398.8837582582582u,0 2399.8602982982984u,0 2399.8612982982986u,1.5 2430.1640395395393u,1.5 2430.1650395395395u,0 2431.1415795795797u,0 2431.14257957958u,1.5 2433.0966596596595u,1.5 2433.0976596596597u,0 2434.0741996996994u,0 2434.0751996996996u,1.5 2436.0292797797797u,1.5 2436.03027977978u,0 2437.0068198198196u,0 2437.00781981982u,1.5 2438.9618998999u,1.5 2438.9628998999u,0 2563.109484984985u,0 2563.1104849849853u,1.5 2564.0870250250246u,1.5 2564.0880250250248u,0 2566.042105105105u,0 2566.043105105105u,1.5 2568.974725225225u,1.5 2568.9757252252252u,0 2569.952265265265u,0 2569.953265265265u,1.5 2570.9298053053053u,1.5 2570.9308053053055u,0 2571.907345345345u,0 2571.9083453453454u,1.5 2601.2335465465467u,1.5 2601.234546546547u,0 2602.2110865865866u,0 2602.212086586587u,1.5 2603.1886266266265u,1.5 2603.1896266266267u,0 2604.1661666666664u,0 2604.1671666666666u,1.5 2605.1437067067063u,1.5 2605.1447067067065u,0 2606.1212467467467u,0 2606.122246746747u,1.5 2607.0987867867866u,1.5 2607.099786786787u,0 2636.424987987988u,0 2636.4259879879883u,1.5 2638.380068068068u,1.5 2638.381068068068u,0 2639.357608108108u,0 2639.358608108108u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2686.27953003003u,0 2686.28053003003u,1.5 2687.25707007007u,1.5 2687.25807007007u,0 2688.2346101101098u,0 2688.23561011011u,1.5 2707.7854109109107u,1.5 2707.786410910911u,0 2708.7629509509507u,0 2708.763950950951u,1.5 2709.740490990991u,1.5 2709.741490990991u,0 2726.3586716716713u,0 2726.3596716716715u,1.5 2727.3362117117117u,1.5 2727.337211711712u,0 2728.3137517517516u,0 2728.314751751752u,1.5 2729.2912917917915u,1.5 2729.2922917917917u,0 2731.2463718718714u,0 2731.2473718718716u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2768.3928933933935u,0 2768.3938933933937u,1.5 2769.3704334334334u,1.5 2769.3714334334336u,0 2770.3479734734733u,0 2770.3489734734735u,1.5 2771.325513513513u,1.5 2771.3265135135134u,0 2772.3030535535536u,0 2772.304053553554u,1.5 2790.876314314314u,1.5 2790.8773143143144u,0 2791.853854354354u,0 2791.8548543543543u,1.5 2792.8313943943945u,1.5 2792.8323943943947u,0 2793.8089344344344u,0 2793.8099344344346u,1.5 2794.7864744744743u,1.5 2794.7874744744745u,0 2814.337275275275u,0 2814.338275275275u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2861.259197197197u,0 2861.260197197197u,1.5 2862.2367372372373u,1.5 2862.2377372372375u,0 2864.191817317317u,0 2864.1928173173173u,1.5 2889.607858358358u,1.5 2889.6088583583582u,0 2890.5853983983984u,0 2890.5863983983986u,1.5 2892.5404784784787u,1.5 2892.541478478479u,0 2893.518018518518u,0 2893.5190185185184u,1.5 2894.4955585585585u,1.5 2894.4965585585587u,0 2897.4281786786787u,0 2897.429178678679u,1.5 2898.4057187187186u,1.5 2898.406718718719u,0 2928.70945995996u,0 2928.71045995996u,1.5 2929.687u,1.5 2929.688u,0 2933.59716016016u,0 2933.59816016016u,1.5 2934.5747002002u,1.5 2934.5757002002u,0 2935.5522402402403u,0 2935.5532402402405u,1.5 2936.52978028028u,1.5 2936.5307802802804u,0 2937.50732032032u,0 2937.5083203203203u,1.5 2939.4624004004004u,1.5 2939.4634004004006u,0 2940.4399404404403u,0 2940.4409404404405u,1.5 2942.39502052052u,1.5 2942.3960205205203u,0 2943.3725605605605u,0 2943.3735605605607u,1.5 3060.677365365365u,1.5 3060.678365365365u,0 3061.6549054054053u,0 3061.6559054054055u,1.5 3063.6099854854856u,1.5 3063.610985485486u,0 3064.587525525525u,0 3064.5885255255253u,1.5 3065.5650655655654u,1.5 3065.5660655655656u,0 3069.4752257257255u,0 3069.4762257257257u,1.5 3070.4527657657654u,1.5 3070.4537657657656u,0 3074.3629259259255u,0 3074.3639259259257u,1.5 3075.340465965966u,1.5 3075.341465965966u,0 3098.8014269269265u,0 3098.8024269269267u,1.5 3099.778966966967u,1.5 3099.779966966967u,0 3102.711587087087u,0 3102.7125870870873u,1.5 3103.689127127127u,1.5 3103.690127127127u,0 3105.644207207207u,0 3105.645207207207u,1.5 3106.621747247247u,1.5 3106.6227472472474u,0 3107.599287287287u,0 3107.6002872872873u,1.5 3108.576827327327u,1.5 3108.577827327327u,0 3109.554367367367u,0 3109.555367367367u,1.5 3132.037788288288u,1.5 3132.0387882882883u,0 3133.0153283283285u,0 3133.0163283283287u,1.5 3134.9704084084083u,1.5 3134.9714084084085u,0 3136.9254884884886u,0 3136.9264884884888u,1.5 3137.9030285285285u,1.5 3137.9040285285287u,0 3161.3639894894895u,0 3161.3649894894897u,1.5 3162.3415295295295u,1.5 3162.3425295295297u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3164.2966096096093u,1.5 3164.2976096096095u,0 3165.2741496496496u,0 3165.27514964965u,1.5 3183.8474104104102u,1.5 3183.8484104104105u,0 3184.82495045045u,0 3184.8259504504504u,1.5 3185.8024904904905u,1.5 3185.8034904904907u,0 3186.7800305305304u,0 3186.7810305305306u,1.5 3187.7575705705704u,1.5 3187.7585705705706u,0 3209.263451451451u,0 3209.2644514514514u,1.5 3229.7917922922925u,1.5 3229.7927922922927u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3269.870933933934u,1.5 3269.871933933934u,0 3270.848473973974u,0 3270.849473973974u,1.5 3271.8260140140137u,1.5 3271.827014014014u,0 3272.803554054054u,0 3272.8045540540543u,1.5 3273.781094094094u,1.5 3273.782094094094u,0 3291.3768148148147u,0 3291.377814814815u,1.5 3312.8826956956955u,1.5 3312.8836956956957u,0 3314.8377757757753u,0 3314.8387757757755u,1.5 3315.8153158158157u,1.5 3315.816315815816u,0 3317.770395895896u,0 3317.771395895896u,1.5 3318.747935935936u,1.5 3318.748935935936u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3337.3211966966965u,1.5 3337.3221966966967u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3361.7596976976974u,1.5 3361.7606976976977u,0 3363.7147777777773u,0 3363.7157777777775u,1.5 3364.6923178178176u,1.5 3364.693317817818u,0 3388.1532787787787u,0 3388.154278778779u,1.5 3389.1308188188186u,1.5 3389.131818818819u,0 3393.040978978979u,0 3393.0419789789794u,1.5 3394.0185190190186u,1.5 3394.019519019019u,0 3394.996059059059u,0 3394.997059059059u,1.5 3398.906219219219u,1.5 3398.9072192192193u,0 3399.883759259259u,0 3399.884759259259u,1.5 3433.12012062062u,1.5 3433.1211206206203u,0 3435.0752007007004u,0 3435.0762007007006u,1.5 3437.0302807807807u,1.5 3437.031280780781u,0 3438.0078208208206u,0 3438.008820820821u,1.5 3438.9853608608605u,1.5 3438.9863608608607u,0 3561.1778658658654u,0 3561.1788658658656u,1.5 3562.155405905906u,1.5 3562.156405905906u,0 3564.110485985986u,0 3564.1114859859863u,1.5 3565.0880260260255u,1.5 3565.0890260260257u,0 3566.065566066066u,0 3566.066566066066u,1.5 3568.998186186186u,1.5 3568.9991861861863u,0 3569.975726226226u,0 3569.976726226226u,1.5 3606.1447077077073u,1.5 3606.1457077077075u,0 3608.0997877877876u,0 3608.100787787788u,1.5 3609.0773278278275u,1.5 3609.0783278278277u,0 3636.4484489489487u,0 3636.449448948949u,1.5 3638.403529029029u,1.5 3638.404529029029u,0 3639.381069069069u,0 3639.382069069069u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3681.4152907907906u,0 3681.4162907907908u,1.5 3682.392830830831u,1.5 3682.393830830831u,0 3685.3254509509507u,0 3685.326450950951u,1.5 3686.302990990991u,1.5 3686.303990990991u,0 3687.280531031031u,0 3687.281531031031u,1.5 3704.8762517517516u,1.5 3704.877251751752u,0 3705.8537917917915u,0 3705.8547917917917u,1.5 3707.8088718718714u,1.5 3707.8098718718716u,0 3708.7864119119117u,0 3708.787411911912u,1.5 3709.7639519519516u,1.5 3709.764951951952u,0 3728.3372127127127u,0 3728.338212712713u,1.5 3729.3147527527526u,1.5 3729.315752752753u,0 3730.292292792793u,0 3730.293292792793u,1.5 3733.2249129129127u,1.5 3733.225912912913u,0 3734.2024529529526u,0 3734.203452952953u,1.5 3746.9104734734733u,1.5 3746.9114734734735u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3770.3714344344344u,0 3770.3724344344346u,1.5 3790.899775275275u,1.5 3790.900775275275u,0 3791.877315315315u,0 3791.8783153153154u,1.5 3792.854855355355u,1.5 3792.8558553553553u,0 3815.338276276276u,0 3815.339276276276u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3862.260198198198u,0 3862.261198198198u,1.5 3864.2152782782778u,1.5 3864.216278278278u,0 3865.192818318318u,0 3865.1938183183183u,1.5 3889.631319319319u,1.5 3889.6323193193193u,0 3890.608859359359u,0 3890.6098593593592u,1.5 3892.5639394394393u,1.5 3892.5649394394395u,0 3893.5414794794797u,0 3893.54247947948u,1.5 3894.519019519519u,1.5 3894.5200195195193u,0 3929.710460960961u,0 3929.711460960961u,1.5 3930.688001001001u,1.5 3930.689001001001u,0 3931.665541041041u,0 3931.666541041041u,1.5 3932.643081081081u,1.5 3932.6440810810814u,0 3934.5981611611614u,0 3934.5991611611616u,1.5 3935.575701201201u,1.5 3935.576701201201u,0 3937.530781281281u,0 3937.5317812812814u,1.5 4064.6109864864866u,1.5 4064.611986486487u,0 4068.5211466466462u,0 4068.5221466466464u,1.5 4069.4986866866866u,1.5 4069.499686686687u,0 4070.4762267267265u,0 4070.4772267267267u,1.5 4071.453766766767u,1.5 4071.454766766767u,0 4103.7125880880885u,0 4103.713588088089u,1.5 4104.690128128128u,1.5 4104.691128128128u,0 4106.645208208208u,0 4106.646208208208u,1.5 4131.083709209209u,1.5 4131.084709209209u,0 4132.061249249249u,0 4132.062249249249u,1.5 4136.948949449449u,1.5 4136.949949449449u,0 4138.904029529529u,0 4138.905029529529u,1.5 4139.881569569569u,1.5 4139.88256956957u,0 4160.40991041041u,0 4160.41091041041u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4162.3649904904905u,0 4162.365990490491u,1.5 4164.32007057057u,1.5 4164.321070570571u,0 4165.297610610611u,0 4165.298610610611u,1.5 4185.825951451451u,1.5 4185.826951451451u,0 4186.8034914914915u,0 4186.804491491492u,1.5 4187.781031531531u,1.5 4187.782031531531u,0 4206.3542922922925u,0 4206.355292292293u,1.5 4207.331832332332u,1.5 4207.332832332332u,0 4208.309372372372u,0 4208.3103723723725u,1.5 4210.264452452452u,1.5 4210.265452452452u,0 4211.2419924924925u,0 4211.242992492493u,1.5 4228.837713213213u,1.5 4228.838713213213u,0 4230.7927932932935u,0 4230.793793293294u,1.5 4231.770333333333u,1.5 4231.771333333333u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4266.961774774775u,1.5 4266.962774774775u,0 4267.939314814815u,0 4267.940314814815u,1.5 4271.849474974975u,1.5 4271.850474974975u,0 4293.355355855856u,0 4293.356355855856u,1.5 4315.838776776777u,1.5 4315.839776776777u,0 4316.816316816817u,0 4316.817316816817u,1.5 4317.793856856857u,1.5 4317.794856856857u,0 4334.412037537537u,0 4334.413037537537u,1.5 4335.389577577577u,1.5 4335.3905775775775u,0 4338.322197697697u,0 4338.323197697698u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4360.805618618619u,1.5 4360.806618618619u,0 4361.783158658659u,0 4361.784158658659u,1.5 4363.738238738738u,1.5 4363.739238738738u,0 4365.693318818819u,0 4365.694318818819u,1.5 4366.670858858859u,1.5 4366.671858858859u,0 4392.086899899899u,0 4392.0878998999u,1.5 4393.06443993994u,1.5 4393.06543993994u,0 4394.04197997998u,0 4394.04297997998u,1.5 4395.01952002002u,1.5 4395.02052002002u,0 4396.9746001001u,0 4396.975600100101u,1.5 4430.210961461462u,1.5 4430.211961461462u,0 4431.188501501501u,0 4431.189501501502u,1.5 4432.166041541541u,1.5 4432.167041541541u,0 4434.121121621622u,0 4434.122121621622u,1.5 4435.098661661662u,1.5 4435.099661661662u,0 4436.076201701701u,0 4436.077201701702u,1.5 4437.053741741741u,1.5 4437.054741741741u,0 4439.008821821822u,0 4439.009821821822u,1.5 4439.986361861862u,1.5 4439.987361861862u,0 4440.963901901901u,0 4440.964901901902u,1.5 4441.941441941942u,1.5 4441.942441941942u,0 4562.178866866867u,0 4562.179866866867u,1.5 4563.156406906906u,1.5 4563.1574069069065u,0 4565.111486986987u,0 4565.112486986987u,1.5 4569.021647147147u,1.5 4569.022647147147u,0 4569.999187187187u,0 4570.000187187187u,1.5 4603.235548548548u,1.5 4603.236548548548u,0 4604.213088588589u,0 4604.214088588589u,1.5 4606.168168668669u,1.5 4606.169168668669u,0 4607.145708708708u,0 4607.1467087087085u,1.5 4608.123248748749u,1.5 4608.124248748749u,0 4634.5168298298295u,0 4634.51782982983u,1.5 4635.49436986987u,1.5 4635.49536986987u,0 4637.44944994995u,0 4637.45044994995u,1.5 4640.38207007007u,1.5 4640.38307007007u,0 4641.35961011011u,0 4641.36061011011u,1.5 4659.932870870871u,1.5 4659.933870870871u,0 4660.91041091091u,0 4660.9114109109105u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4666.775651151151u,0 4666.776651151151u,1.5 4667.753191191191u,1.5 4667.754191191191u,0 4685.348911911911u,0 4685.3499119119115u,1.5 4686.326451951952u,1.5 4686.327451951952u,0 4687.303991991992u,0 4687.304991991992u,1.5 4688.2815320320315u,1.5 4688.282532032032u,0 4689.259072072072u,0 4689.260072072072u,1.5 4705.877252752753u,1.5 4705.878252752753u,0 4706.854792792793u,0 4706.855792792793u,1.5 4707.832332832832u,1.5 4707.833332832833u,0 4708.809872872873u,0 4708.810872872873u,1.5 4709.787412912912u,1.5 4709.7884129129125u,0 4726.405593593594u,0 4726.406593593594u,1.5 4727.383133633633u,1.5 4727.384133633634u,0 4729.338213713713u,0 4729.339213713713u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4770.394895395395u,0 4770.395895395395u,1.5 4772.349975475476u,1.5 4772.350975475476u,0 4773.327515515515u,0 4773.328515515515u,1.5 4792.878316316316u,1.5 4792.879316316316u,0 4795.810936436436u,0 4795.811936436437u,1.5 4796.788476476477u,1.5 4796.789476476477u,0 4815.361737237236u,0 4815.362737237237u,1.5 4816.339277277278u,1.5 4816.340277277278u,0 4817.316817317317u,0 4817.317817317317u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4865.21627927928u,0 4865.21727927928u,1.5 4893.56494044044u,1.5 4893.5659404404405u,0 4895.52002052052u,0 4895.52102052052u,1.5 4896.4975605605605u,1.5 4896.498560560561u,0 4930.711461961962u,0 4930.712461961963u,1.5 4931.689002002002u,1.5 4931.690002002002u,0 4933.644082082082u,0 4933.645082082082u,1.5 4934.621622122122u,1.5 4934.622622122122u,0 4935.599162162162u,0 4935.600162162163u,1.5 4936.576702202202u,1.5 4936.577702202202u,0 4937.554242242241u,0 4937.555242242242u,1.5 4939.509322322322u,1.5 4939.510322322322u,0 4940.486862362362u,0 4940.487862362363u,1.5 5055.8365870870875u,1.5 5055.837587087088u,0 5056.814127127127u,0 5056.815127127127u,1.5 5059.746747247247u,1.5 5059.747747247247u,0 5060.724287287288u,0 5060.725287287288u,1.5 5061.701827327327u,1.5 5061.702827327327u,0 5062.679367367367u,0 5062.680367367368u,1.5 5063.656907407407u,1.5 5063.657907407407u,0 5065.611987487488u,0 5065.612987487488u,1.5 5066.589527527527u,1.5 5066.590527527527u,0 5067.567067567567u,0 5067.568067567568u,1.5 5068.544607607608u,1.5 5068.545607607608u,0 5071.477227727727u,0 5071.478227727727u,1.5 5072.454767767768u,1.5 5072.4557677677685u,0 5103.736049049048u,0 5103.737049049048u,1.5 5105.691129129129u,1.5 5105.692129129129u,0 5106.668669169169u,0 5106.6696691691695u,1.5 5107.646209209209u,1.5 5107.647209209209u,0 5108.623749249249u,0 5108.624749249249u,1.5 5134.0397902902905u,1.5 5134.040790290291u,0 5135.01733033033u,0 5135.01833033033u,1.5 5136.97241041041u,1.5 5136.97341041041u,0 5137.94995045045u,0 5137.95095045045u,1.5 5138.9274904904905u,1.5 5138.928490490491u,0 5161.410911411411u,0 5161.411911411411u,1.5 5163.3659914914915u,1.5 5163.366991491492u,0 5164.343531531531u,0 5164.344531531531u,1.5 5181.939252252252u,1.5 5181.940252252252u,0 5182.9167922922925u,0 5182.917792292293u,1.5 5185.849412412412u,1.5 5185.850412412412u,0 5186.826952452452u,0 5186.827952452452u,1.5 5187.8044924924925u,1.5 5187.805492492493u,0 5207.3552932932935u,0 5207.356293293294u,1.5 5208.332833333333u,1.5 5208.333833333333u,0 5209.310373373373u,0 5209.3113733733735u,1.5 5210.287913413413u,1.5 5210.288913413413u,0 5211.265453453453u,0 5211.266453453453u,1.5 5228.861174174174u,1.5 5228.8621741741745u,0 5230.816254254254u,0 5230.817254254254u,1.5 5231.7937942942945u,1.5 5231.794794294295u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5271.872935935936u,1.5 5271.873935935936u,0 5274.805556056056u,0 5274.806556056056u,1.5 5275.783096096096u,1.5 5275.784096096097u,0 5287.513576576576u,0 5287.5145765765765u,1.5 5288.491116616617u,1.5 5288.492116616617u,0 5292.401276776777u,0 5292.402276776777u,1.5 5313.907157657658u,1.5 5313.908157657658u,0 5315.862237737737u,0 5315.863237737737u,1.5 5316.839777777778u,1.5 5316.840777777778u,0 5339.323198698698u,0 5339.324198698699u,1.5 5359.851539539539u,1.5 5359.852539539539u,0 5360.829079579579u,0 5360.830079579579u,1.5 5365.71677977978u,1.5 5365.71777977978u,0 5392.110360860861u,0 5392.111360860861u,1.5 5393.0879009009u,1.5 5393.088900900901u,0 5396.020521021021u,0 5396.021521021021u,1.5 5433.167042542542u,1.5 5433.168042542542u,0 5434.144582582582u,0 5434.145582582582u,1.5 5435.122122622623u,1.5 5435.123122622623u,0 5436.099662662663u,0 5436.100662662663u,1.5 5437.077202702702u,1.5 5437.078202702703u,0 5442.942442942943u,0 5442.943442942943u,1.5 5443.919982982983u,1.5 5443.920982982983u,0 5557.3146276276275u,0 5557.315627627628u,1.5 5558.292167667668u,1.5 5558.293167667668u,0 5564.157407907907u,0 5564.1584079079075u,1.5 5568.067568068068u,1.5 5568.068568068068u,0 5569.045108108108u,0 5569.0461081081085u,1.5 5601.303929429429u,1.5 5601.30492942943u,0 5602.28146946947u,0 5602.28246946947u,1.5 5604.236549549549u,1.5 5604.237549549549u,0 5606.1916296296295u,0 5606.19262962963u,1.5 5607.16916966967u,1.5 5607.17016966967u,0 5637.47291091091u,0 5637.4739109109105u,1.5 5659.956331831831u,1.5 5659.957331831832u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5662.888951951952u,1.5 5662.889951951952u,0 5685.372372872873u,0 5685.373372872873u,1.5 5686.349912912912u,1.5 5686.3509129129125u,0 5687.327452952953u,0 5687.328452952953u,1.5 5706.878253753754u,1.5 5706.879253753754u,0 5707.855793793794u,0 5707.856793793794u,1.5 5708.833333833833u,1.5 5708.834333833834u,0 5728.384134634634u,0 5728.385134634635u,1.5 5729.361674674675u,1.5 5729.362674674675u,0 5730.339214714714u,0 5730.340214714714u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5769.440816316316u,0 5769.441816316316u,1.5 5770.4183563563565u,1.5 5770.419356356357u,0 5771.395896396396u,0 5771.396896396396u,1.5 5791.924237237236u,1.5 5791.925237237237u,0 5794.8568573573575u,0 5794.857857357358u,1.5 5795.834397397397u,1.5 5795.835397397397u,0 5811.475038038037u,0 5811.476038038038u,1.5 5812.452578078078u,1.5 5812.453578078078u,0 5814.4076581581585u,0 5814.408658158159u,1.5 5816.362738238237u,1.5 5816.363738238238u,0 5817.340278278279u,0 5817.341278278279u,1.5 5833.958458958959u,1.5 5833.95945895896u,0 5834.935998998999u,0 5834.936998998999u,1.5 5836.891079079079u,1.5 5836.892079079079u,0 5837.868619119119u,0 5837.869619119119u,1.5 5839.823699199199u,1.5 5839.824699199199u,0 5861.32958008008u,0 5861.33058008008u,1.5 5862.30712012012u,1.5 5862.30812012012u,0 5863.2846601601605u,0 5863.285660160161u,1.5 5864.2622002002u,1.5 5864.2632002002u,0 5865.239740240239u,0 5865.24074024024u,1.5 5866.217280280281u,1.5 5866.218280280281u,0 5867.19482032032u,0 5867.19582032032u,1.5 5891.633321321321u,1.5 5891.634321321321u,0 5892.6108613613615u,0 5892.611861361362u,1.5 5894.565941441441u,1.5 5894.5669414414415u,0 5896.521021521521u,0 5896.522021521521u,1.5 5897.4985615615615u,1.5 5897.499561561562u,0 5930.734922922923u,0 5930.735922922923u,1.5 5931.712462962963u,1.5 5931.713462962964u,0 5935.622623123123u,0 5935.623623123123u,1.5 5942.465403403403u,1.5 5942.466403403403u,0 5943.442943443443u,0 5943.4439434434435u,1.5 6061.7252882882885u,1.5 6061.726288288289u,0 6063.680368368368u,0 6063.681368368369u,1.5 6064.657908408408u,1.5 6064.658908408408u,0 6065.635448448448u,0 6065.636448448448u,1.5 6066.612988488489u,1.5 6066.613988488489u,0 6074.433308808809u,0 6074.434308808809u,1.5 6075.410848848848u,1.5 6075.411848848848u,0 6103.75951001001u,0 6103.76051001001u,1.5 6104.737050050049u,1.5 6104.738050050049u,0 6105.7145900900905u,0 6105.715590090091u,1.5 6133.085711211211u,1.5 6133.086711211211u,0 6134.063251251251u,0 6134.064251251251u,1.5 6136.995871371371u,1.5 6136.9968713713715u,0 6160.456832332332u,0 6160.457832332332u,1.5 6161.434372372372u,1.5 6161.4353723723725u,0 6162.411912412412u,0 6162.412912412412u,1.5 6163.389452452452u,1.5 6163.390452452452u,0 6164.3669924924925u,0 6164.367992492493u,1.5 6186.850413413413u,1.5 6186.851413413413u,0 6207.378754254254u,0 6207.379754254254u,1.5 6229.862175175175u,1.5 6229.8631751751755u,0 6230.839715215215u,0 6230.840715215215u,1.5 6231.817255255255u,1.5 6231.818255255255u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6251.368056056055u,1.5 6251.369056056055u,0 6252.345596096096u,0 6252.346596096097u,1.5 6267.0086966966965u,1.5 6267.009696696697u,0 6267.986236736736u,0 6267.987236736736u,1.5 6271.8963968968965u,1.5 6271.897396896897u,0 6289.492117617618u,0 6289.493117617618u,1.5 6290.469657657658u,1.5 6290.470657657658u,0 6293.402277777778u,0 6293.403277777778u,1.5 6315.885698698698u,1.5 6315.886698698699u,0 6338.36911961962u,0 6338.37011961962u,1.5 6361.83008058058u,1.5 6361.83108058058u,0 6362.807620620621u,0 6362.808620620621u,1.5 6364.7627007007u,1.5 6364.763700700701u,0 6367.695320820821u,0 6367.696320820821u,1.5 6368.672860860861u,1.5 6368.673860860861u,0 6390.178741741741u,0 6390.179741741741u,1.5 6391.156281781782u,1.5 6391.157281781782u,0 6393.111361861862u,0 6393.112361861862u,1.5 6394.088901901901u,1.5 6394.089901901902u,0 6395.066441941942u,0 6395.067441941942u,1.5 6396.043981981982u,1.5 6396.044981981982u,0 6397.021522022022u,0 6397.022522022022u,1.5 6427.325263263264u,1.5 6427.326263263264u,0 6428.302803303303u,0 6428.3038033033035u,1.5 6432.212963463464u,1.5 6432.213963463464u,0 6433.190503503503u,0 6433.191503503504u,1.5 6434.168043543543u,1.5 6434.169043543543u,0 6435.145583583583u,0 6435.146583583583u,1.5 6436.1231236236235u,1.5 6436.124123623624u,0 6438.078203703703u,0 6438.079203703704u,1.5 6439.055743743743u,1.5 6439.056743743743u,0 6442.965903903903u,0 6442.966903903904u,1.5 6443.943443943944u,1.5 6443.944443943944u,0 6557.338088588589u,0 6557.339088588589u,1.5 6558.3156286286285u,1.5 6558.316628628629u,0 6560.270708708708u,0 6560.2717087087085u,1.5 6561.248248748749u,1.5 6561.249248748749u,0 6562.225788788789u,0 6562.226788788789u,1.5 6563.2033288288285u,1.5 6563.204328828829u,0 6564.180868868869u,0 6564.181868868869u,1.5 6566.135948948949u,1.5 6566.136948948949u,0 6567.113488988989u,0 6567.114488988989u,1.5 6571.023649149149u,1.5 6571.024649149149u,0 6572.001189189189u,0 6572.002189189189u,1.5 6602.30493043043u,1.5 6602.305930430431u,0 6603.282470470471u,0 6603.283470470471u,1.5 6606.215090590591u,1.5 6606.216090590591u,0 6608.170170670671u,0 6608.171170670671u,1.5 6609.14771071071u,1.5 6609.1487107107105u,0 6632.608671671672u,0 6632.609671671672u,1.5 6633.586211711711u,1.5 6633.5872117117115u,0 6634.563751751752u,0 6634.564751751752u,1.5 6635.541291791792u,1.5 6635.542291791792u,0 6636.518831831831u,0 6636.519831831832u,1.5 6640.428991991992u,1.5 6640.429991991992u,0 6641.4065320320315u,0 6641.407532032032u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6684.418293793794u,0 6684.419293793794u,1.5 6685.395833833833u,1.5 6685.396833833834u,0 6687.350913913913u,0 6687.351913913913u,1.5 6707.879254754755u,1.5 6707.880254754755u,0 6725.474975475476u,0 6725.475975475476u,1.5 6726.452515515515u,1.5 6726.453515515515u,0 6729.385135635635u,0 6729.386135635636u,1.5 6730.362675675676u,1.5 6730.363675675676u,0 6731.340215715715u,0 6731.341215715715u,1.5 6747.958396396396u,1.5 6747.959396396396u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6770.441817317317u,0 6770.442817317317u,1.5 6772.396897397397u,1.5 6772.397897397397u,0 6773.374437437437u,0 6773.3754374374375u,1.5 6792.925238238237u,1.5 6792.926238238238u,0 6812.476039039038u,0 6812.477039039039u,1.5 6813.453579079079u,1.5 6813.454579079079u,0 6816.386199199199u,0 6816.387199199199u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6864.285661161161u,0 6864.286661161162u,1.5 6865.263201201201u,1.5 6865.264201201201u,0 6866.24074124124u,0 6866.241741241241u,1.5 6891.656782282283u,1.5 6891.657782282283u,0 6892.634322322322u,0 6892.635322322322u,1.5 6894.589402402402u,1.5 6894.590402402402u,0 6895.566942442442u,0 6895.5679424424425u,1.5 6896.544482482483u,1.5 6896.545482482483u,0 6929.780843843843u,0 6929.7818438438435u,1.5 6930.758383883884u,1.5 6930.759383883884u,0 6935.646084084084u,0 6935.647084084084u,1.5 6937.601164164164u,1.5 6937.602164164165u,0 6938.578704204204u,0 6938.579704204204u,1.5 6943.466404404404u,1.5 6943.467404404404u,0 6944.443944444444u,0 6944.444944444444u,1.5
vbb24 bb24 0 pwl 0,1.5  107.5289044044044u,1.5 107.5299044044044u,0 163.2486866866867u,0 163.2496866866867u,1.5 208.21552852852852u,1.5 208.2165285285285u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 291.3064319319319u,1.5 291.3074319319319u,0 292.28397197197194u,0 292.2849719719719u,1.5 294.23905205205205u,1.5 294.240052052052u,0 334.31819369369373u,0 334.3191936936937u,1.5 335.2957337337337u,1.5 335.2967337337337u,0 337.2508138138138u,0 337.2518138138138u,1.5 391.99305605605605u,1.5 391.994056056056u,0 392.9705960960961u,0 392.97159609609605u,1.5 394.9256761761762u,1.5 394.92667617617616u,0 396.8807562562563u,0 396.88175625625627u,1.5 397.85829629629626u,1.5 397.85929629629624u,0 605.0967847847849u,0 605.0977847847848u,1.5 607.0518648648649u,1.5 607.0528648648649u,0 608.0294049049048u,0 608.0304049049048u,1.5 661.7941071071072u,1.5 661.7951071071071u,0 664.7267272272272u,0 664.7277272272272u,1.5 665.7042672672673u,1.5 665.7052672672672u,0 704.8058688688689u,0 704.8068688688688u,1.5 705.783408908909u,1.5 705.784408908909u,0 708.716029029029u,0 708.7170290290289u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 791.8069324324325u,0 791.8079324324325u,1.5 834.8186941941941u,1.5 834.8196941941941u,0 835.7962342342342u,0 835.7972342342342u,1.5 836.7737742742743u,1.5 836.7747742742743u,0 837.7513143143143u,0 837.7523143143143u,1.5 838.7288543543543u,1.5 838.7298543543543u,0 839.7063943943944u,0 839.7073943943943u,1.5 840.6839344344345u,1.5 840.6849344344345u,0 895.4261766766766u,0 895.4271766766766u,1.5 1106.5748253253253u,1.5 1106.5758253253255u,0 1162.2946076076075u,0 1162.2956076076077u,1.5 1207.2614494494494u,1.5 1207.2624494494496u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1289.3748128128127u,1.5 1289.375812812813u,0 1290.3523528528526u,0 1290.3533528528528u,1.5 1293.2849729729728u,1.5 1293.285972972973u,0 1294.2625130130127u,0 1294.263513013013u,1.5 1295.2400530530529u,1.5 1295.241053053053u,0 1336.2967347347346u,0 1336.2977347347348u,1.5 1337.2742747747748u,1.5 1337.275274774775u,0 1338.251814814815u,0 1338.252814814815u,1.5 1340.2068948948947u,1.5 1340.207894894895u,0 1341.1844349349346u,0 1341.1854349349348u,1.5 1391.0389769769768u,1.5 1391.039976976977u,0 1392.016517017017u,0 1392.017517017017u,1.5 1392.9940570570568u,1.5 1392.995057057057u,0 1393.971597097097u,0 1393.9725970970972u,1.5 1394.9491371371369u,1.5 1394.950137137137u,0 1395.926677177177u,0 1395.9276771771772u,1.5 1396.9042172172171u,1.5 1396.9052172172173u,0 1601.2100855855854u,0 1601.2110855855856u,1.5 1602.1876256256255u,1.5 1602.1886256256257u,0 1605.1202457457457u,0 1605.121245745746u,1.5 1606.0977857857856u,1.5 1606.0987857857858u,0 1608.052865865866u,0 1608.053865865866u,1.5 1609.0304059059058u,1.5 1609.031405905906u,0 1610.007945945946u,0 1610.0089459459462u,1.5 1658.884947947948u,1.5 1658.8859479479481u,0 1659.8624879879878u,0 1659.863487987988u,1.5 1663.7726481481482u,1.5 1663.7736481481484u,0 1706.7844099099098u,0 1706.78540990991u,1.5 1707.76194994995u,1.5 1707.76294994995u,0 1708.73948998999u,0 1708.7404899899902u,1.5 1711.67211011011u,1.5 1711.6731101101102u,0 1712.6496501501501u,0 1712.6506501501503u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1791.8303933933933u,0 1791.8313933933935u,1.5 1792.8079334334332u,1.5 1792.8089334334334u,0 1793.7854734734733u,0 1793.7864734734735u,1.5 1834.842155155155u,1.5 1834.8431551551553u,0 1835.8196951951952u,0 1835.8206951951954u,1.5 1836.7972352352351u,1.5 1836.7982352352353u,0 1837.7747752752753u,0 1837.7757752752755u,1.5 1838.7523153153154u,1.5 1838.7533153153156u,0 1887.6293173173174u,0 1887.6303173173176u,1.5 1888.6068573573573u,1.5 1888.6078573573575u,0 1890.5619374374373u,0 1890.5629374374375u,1.5 1891.5394774774772u,1.5 1891.5404774774775u,0 1893.4945575575573u,0 1893.4955575575575u,1.5 1894.4720975975974u,1.5 1894.4730975975976u,0 1895.4496376376374u,0 1895.4506376376376u,1.5 2104.643206206206u,1.5 2104.644206206206u,0 2107.575826326326u,0 2107.576826326326u,1.5 2108.553366366366u,1.5 2108.554366366366u,0 2112.463526526526u,0 2112.4645265265262u,1.5 2113.4410665665664u,1.5 2113.4420665665666u,0 2161.3405285285285u,0 2161.3415285285287u,1.5 2166.228228728729u,1.5 2166.229228728729u,0 2167.2057687687684u,0 2167.2067687687686u,1.5 2206.30737037037u,1.5 2206.30837037037u,0 2207.2849104104102u,0 2207.2859104104105u,1.5 2209.2399904904905u,1.5 2209.2409904904907u,0 2250.296672172172u,0 2250.297672172172u,1.5 2291.3533538538536u,1.5 2291.354353853854u,0 2292.330893893894u,0 2292.331893893894u,1.5 2294.285973973974u,1.5 2294.286973973974u,0 2338.2752757757753u,0 2338.2762757757755u,1.5 2388.1298178178176u,1.5 2388.130817817818u,0 2389.1073578578576u,0 2389.1083578578578u,1.5 2393.0175180180177u,1.5 2393.018518018018u,0 2393.995058058058u,0 2393.996058058058u,1.5 2394.972598098098u,1.5 2394.973598098098u,0 2395.9501381381383u,0 2395.9511381381385u,1.5 2396.927678178178u,1.5 2396.9286781781784u,0 2398.882758258258u,0 2398.8837582582582u,1.5 2399.8602982982984u,1.5 2399.8612982982986u,0 2601.2335465465467u,0 2601.234546546547u,1.5 2602.2110865865866u,1.5 2602.212086586587u,0 2603.1886266266265u,0 2603.1896266266267u,1.5 2604.1661666666664u,1.5 2604.1671666666666u,0 2605.1437067067063u,0 2605.1447067067065u,1.5 2606.1212467467467u,1.5 2606.122246746747u,0 2607.0987867867866u,0 2607.099786786787u,1.5 2660.863488988989u,1.5 2660.8644889889893u,0 2661.841029029029u,0 2661.842029029029u,1.5 2662.818569069069u,1.5 2662.819569069069u,0 2663.796109109109u,0 2663.797109109109u,1.5 2664.773649149149u,1.5 2664.7746491491494u,0 2707.7854109109107u,0 2707.786410910911u,1.5 2708.7629509509507u,1.5 2708.763950950951u,0 2709.740490990991u,0 2709.741490990991u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2790.876314314314u,0 2790.8773143143144u,1.5 2791.853854354354u,1.5 2791.8548543543543u,0 2792.8313943943945u,0 2792.8323943943947u,1.5 2793.8089344344344u,1.5 2793.8099344344346u,0 2794.7864744744743u,0 2794.7874744744745u,1.5 2835.843156156156u,1.5 2835.8441561561563u,0 2836.820696196196u,0 2836.821696196196u,1.5 2838.775776276276u,1.5 2838.776776276276u,0 2889.607858358358u,0 2889.6088583583582u,1.5 2890.5853983983984u,1.5 2890.5863983983986u,0 2892.5404784784787u,0 2892.541478478479u,1.5 2893.518018518518u,1.5 2893.5190185185184u,0 2894.4955585585585u,0 2894.4965585585587u,1.5 2897.4281786786787u,1.5 2897.429178678679u,0 2898.4057187187186u,0 2898.406718718719u,1.5 3098.8014269269265u,1.5 3098.8024269269267u,0 3099.778966966967u,0 3099.779966966967u,1.5 3102.711587087087u,1.5 3102.7125870870873u,0 3103.689127127127u,0 3103.690127127127u,1.5 3105.644207207207u,1.5 3105.645207207207u,0 3106.621747247247u,0 3106.6227472472474u,1.5 3107.599287287287u,1.5 3107.6002872872873u,0 3108.576827327327u,0 3108.577827327327u,1.5 3109.554367367367u,1.5 3109.555367367367u,0 3161.3639894894895u,0 3161.3649894894897u,1.5 3162.3415295295295u,1.5 3162.3425295295297u,0 3163.3190695695694u,0 3163.3200695695696u,1.5 3164.2966096096093u,1.5 3164.2976096096095u,0 3165.2741496496496u,0 3165.27514964965u,1.5 3209.263451451451u,1.5 3209.2644514514514u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3291.3768148148147u,1.5 3291.377814814815u,0 3336.3436566566565u,0 3336.3446566566568u,1.5 3337.3211966966965u,1.5 3337.3221966966967u,0 3339.2762767767763u,0 3339.2772767767765u,1.5 3388.1532787787787u,1.5 3388.154278778779u,0 3389.1308188188186u,0 3389.131818818819u,1.5 3393.040978978979u,1.5 3393.0419789789794u,0 3394.0185190190186u,0 3394.019519019019u,1.5 3394.996059059059u,1.5 3394.997059059059u,0 3398.906219219219u,0 3398.9072192192193u,1.5 3399.883759259259u,1.5 3399.884759259259u,0 3606.1447077077073u,0 3606.1457077077075u,1.5 3608.0997877877876u,1.5 3608.100787787788u,0 3609.0773278278275u,0 3609.0783278278277u,1.5 3660.8869499499497u,1.5 3660.88794994995u,0 3661.86448998999u,0 3661.8654899899902u,1.5 3663.81957007007u,1.5 3663.82057007007u,0 3704.8762517517516u,0 3704.877251751752u,1.5 3705.8537917917915u,1.5 3705.8547917917917u,0 3707.8088718718714u,0 3707.8098718718716u,1.5 3708.7864119119117u,1.5 3708.787411911912u,0 3709.7639519519516u,0 3709.764951951952u,1.5 3746.9104734734733u,1.5 3746.9114734734735u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3790.899775275275u,0 3790.900775275275u,1.5 3791.877315315315u,1.5 3791.8783153153154u,0 3792.854855355355u,0 3792.8558553553553u,1.5 3834.8890770770768u,1.5 3834.890077077077u,0 3835.8666171171167u,0 3835.867617117117u,1.5 3838.7992372372373u,1.5 3838.8002372372375u,0 3889.631319319319u,0 3889.6323193193193u,1.5 3890.608859359359u,1.5 3890.6098593593592u,0 3892.5639394394393u,0 3892.5649394394395u,1.5 3893.5414794794797u,1.5 3893.54247947948u,0 3894.519019519519u,0 3894.5200195195193u,1.5 4103.7125880880885u,1.5 4103.713588088089u,0 4104.690128128128u,0 4104.691128128128u,1.5 4106.645208208208u,1.5 4106.646208208208u,0 4160.40991041041u,0 4160.41091041041u,1.5 4161.38745045045u,1.5 4161.38845045045u,0 4162.3649904904905u,0 4162.365990490491u,1.5 4164.32007057057u,1.5 4164.321070570571u,0 4165.297610610611u,0 4165.298610610611u,1.5 4206.3542922922925u,1.5 4206.355292292293u,0 4207.331832332332u,0 4207.332832332332u,1.5 4208.309372372372u,1.5 4208.3103723723725u,0 4210.264452452452u,0 4210.265452452452u,1.5 4211.2419924924925u,1.5 4211.242992492493u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4293.355355855856u,1.5 4293.356355855856u,0 4334.412037537537u,0 4334.413037537537u,1.5 4335.389577577577u,1.5 4335.3905775775775u,0 4338.322197697697u,0 4338.323197697698u,1.5 4340.277277777778u,1.5 4340.278277777778u,0 4341.254817817818u,0 4341.255817817818u,1.5 4392.086899899899u,1.5 4392.0878998999u,0 4393.06443993994u,0 4393.06543993994u,1.5 4394.04197997998u,1.5 4394.04297997998u,0 4395.01952002002u,0 4395.02052002002u,1.5 4396.9746001001u,1.5 4396.975600100101u,0 4603.235548548548u,0 4603.236548548548u,1.5 4604.213088588589u,1.5 4604.214088588589u,0 4606.168168668669u,0 4606.169168668669u,1.5 4607.145708708708u,1.5 4607.1467087087085u,0 4608.123248748749u,0 4608.124248748749u,1.5 4659.932870870871u,1.5 4659.933870870871u,0 4660.91041091091u,0 4660.9114109109105u,1.5 4661.887950950951u,1.5 4661.888950950951u,0 4663.8430310310305u,0 4663.844031031031u,1.5 4664.820571071071u,1.5 4664.821571071071u,0 4666.775651151151u,0 4666.776651151151u,1.5 4667.753191191191u,1.5 4667.754191191191u,0 4705.877252752753u,0 4705.878252752753u,1.5 4706.854792792793u,1.5 4706.855792792793u,0 4707.832332832832u,0 4707.833332832833u,1.5 4708.809872872873u,1.5 4708.810872872873u,0 4709.787412912912u,0 4709.7884129129125u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4792.878316316316u,0 4792.879316316316u,1.5 4795.810936436436u,1.5 4795.811936436437u,0 4796.788476476477u,0 4796.789476476477u,1.5 4836.867618118118u,1.5 4836.868618118118u,0 4837.8451581581585u,0 4837.846158158159u,1.5 4838.822698198198u,1.5 4838.823698198198u,0 4893.56494044044u,0 4893.5659404404405u,1.5 4895.52002052052u,1.5 4895.52102052052u,0 4896.4975605605605u,0 4896.498560560561u,1.5 5103.736049049048u,1.5 5103.737049049048u,0 5105.691129129129u,0 5105.692129129129u,1.5 5106.668669169169u,1.5 5106.6696691691695u,0 5107.646209209209u,0 5107.647209209209u,1.5 5108.623749249249u,1.5 5108.624749249249u,0 5161.410911411411u,0 5161.411911411411u,1.5 5163.3659914914915u,1.5 5163.366991491492u,0 5164.343531531531u,0 5164.344531531531u,1.5 5207.3552932932935u,1.5 5207.356293293294u,0 5208.332833333333u,0 5208.333833333333u,1.5 5209.310373373373u,1.5 5209.3113733733735u,0 5210.287913413413u,0 5210.288913413413u,1.5 5211.265453453453u,1.5 5211.266453453453u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5287.513576576576u,1.5 5287.5145765765765u,0 5288.491116616617u,0 5288.492116616617u,1.5 5292.401276776777u,1.5 5292.402276776777u,0 5339.323198698698u,0 5339.324198698699u,1.5 5392.110360860861u,1.5 5392.111360860861u,0 5393.0879009009u,0 5393.088900900901u,1.5 5396.020521021021u,1.5 5396.021521021021u,0 5601.303929429429u,0 5601.30492942943u,1.5 5602.28146946947u,1.5 5602.28246946947u,0 5604.236549549549u,0 5604.237549549549u,1.5 5606.1916296296295u,1.5 5606.19262962963u,0 5607.16916966967u,0 5607.17016966967u,1.5 5659.956331831831u,1.5 5659.957331831832u,0 5661.911411911911u,0 5661.9124119119115u,1.5 5662.888951951952u,1.5 5662.889951951952u,0 5706.878253753754u,0 5706.879253753754u,1.5 5707.855793793794u,1.5 5707.856793793794u,0 5708.833333833833u,0 5708.834333833834u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5791.924237237236u,0 5791.925237237237u,1.5 5794.8568573573575u,1.5 5794.857857357358u,0 5795.834397397397u,0 5795.835397397397u,1.5 5833.958458958959u,1.5 5833.95945895896u,0 5834.935998998999u,0 5834.936998998999u,1.5 5836.891079079079u,1.5 5836.892079079079u,0 5837.868619119119u,0 5837.869619119119u,1.5 5839.823699199199u,1.5 5839.824699199199u,0 5891.633321321321u,0 5891.634321321321u,1.5 5892.6108613613615u,1.5 5892.611861361362u,0 5894.565941441441u,0 5894.5669414414415u,1.5 5896.521021521521u,1.5 5896.522021521521u,0 5897.4985615615615u,0 5897.499561561562u,1.5 6103.75951001001u,1.5 6103.76051001001u,0 6104.737050050049u,0 6104.738050050049u,1.5 6105.7145900900905u,1.5 6105.715590090091u,0 6160.456832332332u,0 6160.457832332332u,1.5 6161.434372372372u,1.5 6161.4353723723725u,0 6162.411912412412u,0 6162.412912412412u,1.5 6163.389452452452u,1.5 6163.390452452452u,0 6164.3669924924925u,0 6164.367992492493u,1.5 6207.378754254254u,1.5 6207.379754254254u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6251.368056056055u,1.5 6251.369056056055u,0 6252.345596096096u,0 6252.346596096097u,1.5 6289.492117617618u,1.5 6289.493117617618u,0 6290.469657657658u,0 6290.470657657658u,1.5 6293.402277777778u,1.5 6293.403277777778u,0 6338.36911961962u,0 6338.37011961962u,1.5 6390.178741741741u,1.5 6390.179741741741u,0 6391.156281781782u,0 6391.157281781782u,1.5 6393.111361861862u,1.5 6393.112361861862u,0 6394.088901901901u,0 6394.089901901902u,1.5 6395.066441941942u,1.5 6395.067441941942u,0 6396.043981981982u,0 6396.044981981982u,1.5 6397.021522022022u,1.5 6397.022522022022u,0 6602.30493043043u,0 6602.305930430431u,1.5 6603.282470470471u,1.5 6603.283470470471u,0 6606.215090590591u,0 6606.216090590591u,1.5 6608.170170670671u,1.5 6608.171170670671u,0 6609.14771071071u,0 6609.1487107107105u,1.5 6660.957332832832u,1.5 6660.958332832833u,0 6661.934872872873u,0 6661.935872872873u,1.5 6663.889952952953u,1.5 6663.890952952953u,0 6707.879254754755u,0 6707.880254754755u,1.5 6747.958396396396u,1.5 6747.959396396396u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6792.925238238237u,0 6792.926238238238u,1.5 6837.89208008008u,1.5 6837.89308008008u,0 6891.656782282283u,0 6891.657782282283u,1.5 6892.634322322322u,1.5 6892.635322322322u,0 6894.589402402402u,0 6894.590402402402u,1.5 6895.566942442442u,1.5 6895.5679424424425u,0 6896.544482482483u,0 6896.545482482483u,1.5
vbb25 bb25 0 pwl 0,1.5  163.2486866866867u,1.5 163.2496866866867u,0 249.27221021021023u,0 249.2732102102102u,1.5 250.24975025025026u,1.5 250.25075025025023u,0 251.22729029029028u,0 251.22829029029026u,1.5 334.31819369369373u,1.5 334.3191936936937u,0 335.2957337337337u,0 335.2967337337337u,1.5 337.2508138138138u,1.5 337.2518138138138u,0 661.7941071071072u,0 661.7951071071071u,1.5 664.7267272272272u,1.5 664.7277272272272u,0 665.7042672672673u,0 665.7052672672672u,1.5 749.7727107107107u,1.5 749.7737107107107u,0 750.7502507507508u,0 750.7512507507507u,1.5 751.7277907907908u,1.5 751.7287907907908u,0 834.8186941941941u,0 834.8196941941941u,1.5 835.7962342342342u,1.5 835.7972342342342u,0 836.7737742742743u,0 836.7747742742743u,1.5 837.7513143143143u,1.5 837.7523143143143u,0 838.7288543543543u,0 838.7298543543543u,1.5 839.7063943943944u,1.5 839.7073943943943u,0 840.6839344344345u,0 840.6849344344345u,1.5 1162.2946076076075u,1.5 1162.2956076076077u,0 1250.273211211211u,0 1250.2742112112112u,1.5 1336.2967347347346u,1.5 1336.2977347347348u,0 1337.2742747747748u,0 1337.275274774775u,1.5 1338.251814814815u,1.5 1338.252814814815u,0 1340.2068948948947u,0 1340.207894894895u,1.5 1341.1844349349346u,1.5 1341.1854349349348u,0 1658.884947947948u,0 1658.8859479479481u,1.5 1659.8624879879878u,1.5 1659.863487987988u,0 1663.7726481481482u,0 1663.7736481481484u,1.5 1749.7961716716716u,1.5 1749.7971716716718u,0 1750.7737117117115u,0 1750.7747117117117u,1.5 1751.7512517517516u,1.5 1751.7522517517518u,0 1834.842155155155u,0 1834.8431551551553u,1.5 1835.8196951951952u,1.5 1835.8206951951954u,0 1836.7972352352351u,0 1836.7982352352353u,1.5 1837.7747752752753u,1.5 1837.7757752752755u,0 1838.7523153153154u,0 1838.7533153153156u,1.5 2161.3405285285285u,1.5 2161.3415285285287u,0 2166.228228728729u,0 2166.229228728729u,1.5 2167.2057687687684u,1.5 2167.2067687687686u,0 2250.296672172172u,0 2250.297672172172u,1.5 2338.2752757757753u,1.5 2338.2762757757755u,0 2660.863488988989u,0 2660.8644889889893u,1.5 2661.841029029029u,1.5 2661.842029029029u,0 2662.818569069069u,0 2662.819569069069u,1.5 2663.796109109109u,1.5 2663.797109109109u,0 2664.773649149149u,0 2664.7746491491494u,1.5 2749.819632632633u,1.5 2749.820632632633u,0 2835.843156156156u,0 2835.8441561561563u,1.5 2836.820696196196u,1.5 2836.821696196196u,0 2838.775776276276u,0 2838.776776276276u,1.5 3161.3639894894895u,1.5 3161.3649894894897u,0 3162.3415295295295u,0 3162.3425295295297u,1.5 3163.3190695695694u,1.5 3163.3200695695696u,0 3164.2966096096093u,0 3164.2976096096095u,1.5 3165.2741496496496u,1.5 3165.27514964965u,0 3248.365053053053u,0 3248.3660530530533u,1.5 3249.342593093093u,1.5 3249.343593093093u,0 3251.297673173173u,0 3251.298673173173u,1.5 3252.275213213213u,1.5 3252.2762132132134u,0 3253.252753253253u,0 3253.2537532532533u,1.5 3336.3436566566565u,1.5 3336.3446566566568u,0 3337.3211966966965u,0 3337.3221966966967u,1.5 3339.2762767767763u,1.5 3339.2772767767765u,0 3660.8869499499497u,0 3660.88794994995u,1.5 3661.86448998999u,1.5 3661.8654899899902u,0 3663.81957007007u,0 3663.82057007007u,1.5 3746.9104734734733u,1.5 3746.9114734734735u,0 3747.888013513513u,0 3747.8890135135134u,1.5 3748.8655535535536u,1.5 3748.866553553554u,0 3749.8430935935935u,0 3749.8440935935937u,1.5 3750.820633633634u,1.5 3750.821633633634u,0 3751.7981736736733u,0 3751.7991736736735u,1.5 3752.7757137137137u,1.5 3752.776713713714u,0 3834.8890770770768u,0 3834.890077077077u,1.5 3835.8666171171167u,1.5 3835.867617117117u,0 3838.7992372372373u,0 3838.8002372372375u,1.5 4160.40991041041u,1.5 4160.41091041041u,0 4161.38745045045u,0 4161.38845045045u,1.5 4162.3649904904905u,1.5 4162.365990490491u,0 4164.32007057057u,0 4164.321070570571u,1.5 4165.297610610611u,1.5 4165.298610610611u,0 4249.366054054053u,0 4249.367054054053u,1.5 4250.343594094094u,1.5 4250.344594094095u,0 4251.321134134134u,0 4251.322134134134u,1.5 4334.412037537537u,1.5 4334.413037537537u,0 4335.389577577577u,0 4335.3905775775775u,1.5 4338.322197697697u,1.5 4338.323197697698u,0 4340.277277777778u,0 4340.278277777778u,1.5 4341.254817817818u,1.5 4341.255817817818u,0 4659.932870870871u,0 4659.933870870871u,1.5 4660.91041091091u,1.5 4660.9114109109105u,0 4661.887950950951u,0 4661.888950950951u,1.5 4663.8430310310305u,1.5 4663.844031031031u,0 4664.820571071071u,0 4664.821571071071u,1.5 4666.775651151151u,1.5 4666.776651151151u,0 4667.753191191191u,0 4667.754191191191u,1.5 4747.911474474475u,1.5 4747.912474474475u,0 4748.889014514514u,0 4748.890014514514u,1.5 4749.866554554554u,1.5 4749.867554554554u,0 4751.821634634634u,0 4751.822634634635u,1.5 4752.799174674675u,1.5 4752.800174674675u,0 4836.867618118118u,0 4836.868618118118u,1.5 4837.8451581581585u,1.5 4837.846158158159u,0 4838.822698198198u,0 4838.823698198198u,1.5 5161.410911411411u,1.5 5161.411911411411u,0 5163.3659914914915u,0 5163.366991491492u,1.5 5164.343531531531u,1.5 5164.344531531531u,0 5249.389515015015u,0 5249.390515015015u,1.5 5250.367055055054u,1.5 5250.368055055054u,0 5251.344595095095u,0 5251.345595095096u,1.5 5339.323198698698u,1.5 5339.324198698699u,0 5659.956331831831u,0 5659.957331831832u,1.5 5661.911411911911u,1.5 5661.9124119119115u,0 5662.888951951952u,0 5662.889951951952u,1.5 5750.867555555555u,1.5 5750.868555555555u,0 5833.958458958959u,0 5833.95945895896u,1.5 5834.935998998999u,1.5 5834.936998998999u,0 5836.891079079079u,0 5836.892079079079u,1.5 5837.868619119119u,1.5 5837.869619119119u,0 5839.823699199199u,0 5839.824699199199u,1.5 6160.456832332332u,1.5 6160.457832332332u,0 6161.434372372372u,0 6161.4353723723725u,1.5 6162.411912412412u,1.5 6162.412912412412u,0 6163.389452452452u,0 6163.390452452452u,1.5 6164.3669924924925u,1.5 6164.367992492493u,0 6248.435435935936u,0 6248.436435935936u,1.5 6249.412975975976u,1.5 6249.413975975976u,0 6250.390516016016u,0 6250.391516016016u,1.5 6251.368056056055u,1.5 6251.369056056055u,0 6252.345596096096u,0 6252.346596096097u,1.5 6338.36911961962u,1.5 6338.37011961962u,0 6660.957332832832u,0 6660.958332832833u,1.5 6661.934872872873u,1.5 6661.935872872873u,0 6663.889952952953u,0 6663.890952952953u,1.5 6747.958396396396u,1.5 6747.959396396396u,0 6748.935936436436u,0 6748.936936436437u,1.5 6750.891016516516u,1.5 6750.892016516516u,0 6837.89208008008u,0 6837.89308008008u,1.5
vbb26 bb26 0 pwl 0,1.5  249.27221021021023u,1.5 249.2732102102102u,0 250.24975025025026u,0 250.25075025025023u,1.5 251.22729029029028u,1.5 251.22829029029026u,0 749.7727107107107u,0 749.7737107107107u,1.5 750.7502507507508u,1.5 750.7512507507507u,0 751.7277907907908u,0 751.7287907907908u,1.5 1250.273211211211u,1.5 1250.2742112112112u,0 1749.7961716716716u,0 1749.7971716716718u,1.5 1750.7737117117115u,1.5 1750.7747117117117u,0 1751.7512517517516u,0 1751.7522517517518u,1.5 2250.296672172172u,1.5 2250.297672172172u,0 2749.819632632633u,0 2749.820632632633u,1.5 3248.365053053053u,1.5 3248.3660530530533u,0 3249.342593093093u,0 3249.343593093093u,1.5 3251.297673173173u,1.5 3251.298673173173u,0 3252.275213213213u,0 3252.2762132132134u,1.5 3253.252753253253u,1.5 3253.2537532532533u,0 3746.9104734734733u,0 3746.9114734734735u,1.5 3747.888013513513u,1.5 3747.8890135135134u,0 3748.8655535535536u,0 3748.866553553554u,1.5 3749.8430935935935u,1.5 3749.8440935935937u,0 3750.820633633634u,0 3750.821633633634u,1.5 3751.7981736736733u,1.5 3751.7991736736735u,0 3752.7757137137137u,0 3752.776713713714u,1.5 4249.366054054053u,1.5 4249.367054054053u,0 4250.343594094094u,0 4250.344594094095u,1.5 4251.321134134134u,1.5 4251.322134134134u,0 4747.911474474475u,0 4747.912474474475u,1.5 4748.889014514514u,1.5 4748.890014514514u,0 4749.866554554554u,0 4749.867554554554u,1.5 4751.821634634634u,1.5 4751.822634634635u,0 4752.799174674675u,0 4752.800174674675u,1.5 5249.389515015015u,1.5 5249.390515015015u,0 5250.367055055054u,0 5250.368055055054u,1.5 5251.344595095095u,1.5 5251.345595095096u,0 5750.867555555555u,0 5750.868555555555u,1.5 6248.435435935936u,1.5 6248.436435935936u,0 6249.412975975976u,0 6249.413975975976u,1.5 6250.390516016016u,1.5 6250.391516016016u,0 6251.368056056055u,0 6251.369056056055u,1.5 6252.345596096096u,1.5 6252.346596096097u,0 6747.958396396396u,0 6747.959396396396u,1.5 6748.935936436436u,1.5 6748.936936436437u,0 6750.891016516516u,0 6750.892016516516u,1.5
